VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplier
  CLASS BLOCK ;
  FOREIGN multiplier ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END clk
  PIN input_a1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END input_a1[0]
  PIN input_a1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.370 0.000 928.650 4.000 ;
    END
  END input_a1[10]
  PIN input_a1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 655.560 1000.000 656.160 ;
    END
  END input_a1[11]
  PIN input_a1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 996.000 510.050 1000.000 ;
    END
  END input_a1[12]
  PIN input_a1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 427.080 1000.000 427.680 ;
    END
  END input_a1[13]
  PIN input_a1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 579.400 1000.000 580.000 ;
    END
  END input_a1[14]
  PIN input_a1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 198.600 1000.000 199.200 ;
    END
  END input_a1[15]
  PIN input_a1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 960.200 1000.000 960.800 ;
    END
  END input_a1[1]
  PIN input_a1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 996.000 45.450 1000.000 ;
    END
  END input_a1[2]
  PIN input_a1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 913.960 4.000 914.560 ;
    END
  END input_a1[3]
  PIN input_a1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.850 0.000 877.130 4.000 ;
    END
  END input_a1[4]
  PIN input_a1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 996.000 458.530 1000.000 ;
    END
  END input_a1[5]
  PIN input_a1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 996.000 716.130 1000.000 ;
    END
  END input_a1[6]
  PIN input_a1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END input_a1[7]
  PIN input_a1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 122.440 1000.000 123.040 ;
    END
  END input_a1[8]
  PIN input_a1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 503.240 1000.000 503.840 ;
    END
  END input_a1[9]
  PIN input_b1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END input_b1[0]
  PIN input_b1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END input_b1[10]
  PIN input_b1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 884.040 1000.000 884.640 ;
    END
  END input_b1[11]
  PIN input_b1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 996.000 613.090 1000.000 ;
    END
  END input_b1[12]
  PIN input_b1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END input_b1[13]
  PIN input_b1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.120 4.000 990.720 ;
    END
  END input_b1[14]
  PIN input_b1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END input_b1[15]
  PIN input_b1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END input_b1[1]
  PIN input_b1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END input_b1[2]
  PIN input_b1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END input_b1[3]
  PIN input_b1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 996.000 355.490 1000.000 ;
    END
  END input_b1[4]
  PIN input_b1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END input_b1[5]
  PIN input_b1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 996.000 664.610 1000.000 ;
    END
  END input_b1[6]
  PIN input_b1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 996.000 148.490 1000.000 ;
    END
  END input_b1[7]
  PIN input_b1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 0.000 980.170 4.000 ;
    END
  END input_b1[8]
  PIN input_b1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END input_b1[9]
  PIN product[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 46.280 1000.000 46.880 ;
    END
  END product[0]
  PIN product[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 996.000 819.170 1000.000 ;
    END
  END product[10]
  PIN product[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END product[11]
  PIN product[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 996.000 252.450 1000.000 ;
    END
  END product[12]
  PIN product[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END product[13]
  PIN product[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END product[14]
  PIN product[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 996.000 767.650 1000.000 ;
    END
  END product[15]
  PIN product[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END product[16]
  PIN product[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 807.880 1000.000 808.480 ;
    END
  END product[17]
  PIN product[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 996.000 561.570 1000.000 ;
    END
  END product[18]
  PIN product[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END product[19]
  PIN product[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END product[1]
  PIN product[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 996.000 200.930 1000.000 ;
    END
  END product[20]
  PIN product[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.450 996.000 973.730 1000.000 ;
    END
  END product[21]
  PIN product[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END product[22]
  PIN product[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 731.720 1000.000 732.320 ;
    END
  END product[23]
  PIN product[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END product[24]
  PIN product[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END product[25]
  PIN product[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 274.760 1000.000 275.360 ;
    END
  END product[26]
  PIN product[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END product[27]
  PIN product[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END product[28]
  PIN product[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END product[29]
  PIN product[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END product[2]
  PIN product[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END product[30]
  PIN product[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 996.000 922.210 1000.000 ;
    END
  END product[31]
  PIN product[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 996.000 870.690 1000.000 ;
    END
  END product[3]
  PIN product[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 996.000 303.970 1000.000 ;
    END
  END product[4]
  PIN product[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 996.000 407.010 1000.000 ;
    END
  END product[5]
  PIN product[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END product[6]
  PIN product[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END product[7]
  PIN product[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 996.000 96.970 1000.000 ;
    END
  END product[8]
  PIN product[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 350.920 1000.000 351.520 ;
    END
  END product[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 204.720 10.640 206.320 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.720 10.640 406.320 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.720 10.640 606.320 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 804.720 10.640 806.320 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.720 10.640 106.320 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.720 10.640 306.320 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.720 10.640 506.320 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.720 10.640 706.320 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.720 10.640 906.320 987.600 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.835 987.445 ;
      LAYER met1 ;
        RECT 0.070 9.560 994.895 987.600 ;
      LAYER met2 ;
        RECT 0.100 995.720 44.890 996.000 ;
        RECT 45.730 995.720 96.410 996.000 ;
        RECT 97.250 995.720 147.930 996.000 ;
        RECT 148.770 995.720 200.370 996.000 ;
        RECT 201.210 995.720 251.890 996.000 ;
        RECT 252.730 995.720 303.410 996.000 ;
        RECT 304.250 995.720 354.930 996.000 ;
        RECT 355.770 995.720 406.450 996.000 ;
        RECT 407.290 995.720 457.970 996.000 ;
        RECT 458.810 995.720 509.490 996.000 ;
        RECT 510.330 995.720 561.010 996.000 ;
        RECT 561.850 995.720 612.530 996.000 ;
        RECT 613.370 995.720 664.050 996.000 ;
        RECT 664.890 995.720 715.570 996.000 ;
        RECT 716.410 995.720 767.090 996.000 ;
        RECT 767.930 995.720 818.610 996.000 ;
        RECT 819.450 995.720 870.130 996.000 ;
        RECT 870.970 995.720 921.650 996.000 ;
        RECT 922.490 995.720 973.170 996.000 ;
        RECT 974.010 995.720 989.830 996.000 ;
        RECT 0.100 4.280 989.830 995.720 ;
        RECT 0.650 4.000 51.330 4.280 ;
        RECT 52.170 4.000 102.850 4.280 ;
        RECT 103.690 4.000 154.370 4.280 ;
        RECT 155.210 4.000 205.890 4.280 ;
        RECT 206.730 4.000 257.410 4.280 ;
        RECT 258.250 4.000 308.930 4.280 ;
        RECT 309.770 4.000 360.450 4.280 ;
        RECT 361.290 4.000 411.970 4.280 ;
        RECT 412.810 4.000 463.490 4.280 ;
        RECT 464.330 4.000 515.010 4.280 ;
        RECT 515.850 4.000 566.530 4.280 ;
        RECT 567.370 4.000 618.050 4.280 ;
        RECT 618.890 4.000 669.570 4.280 ;
        RECT 670.410 4.000 721.090 4.280 ;
        RECT 721.930 4.000 772.610 4.280 ;
        RECT 773.450 4.000 824.130 4.280 ;
        RECT 824.970 4.000 876.570 4.280 ;
        RECT 877.410 4.000 928.090 4.280 ;
        RECT 928.930 4.000 979.610 4.280 ;
        RECT 980.450 4.000 989.830 4.280 ;
      LAYER met3 ;
        RECT 4.400 989.720 996.000 990.585 ;
        RECT 4.000 961.200 996.000 989.720 ;
        RECT 4.000 959.800 995.600 961.200 ;
        RECT 4.000 914.960 996.000 959.800 ;
        RECT 4.400 913.560 996.000 914.960 ;
        RECT 4.000 885.040 996.000 913.560 ;
        RECT 4.000 883.640 995.600 885.040 ;
        RECT 4.000 838.800 996.000 883.640 ;
        RECT 4.400 837.400 996.000 838.800 ;
        RECT 4.000 808.880 996.000 837.400 ;
        RECT 4.000 807.480 995.600 808.880 ;
        RECT 4.000 762.640 996.000 807.480 ;
        RECT 4.400 761.240 996.000 762.640 ;
        RECT 4.000 732.720 996.000 761.240 ;
        RECT 4.000 731.320 995.600 732.720 ;
        RECT 4.000 686.480 996.000 731.320 ;
        RECT 4.400 685.080 996.000 686.480 ;
        RECT 4.000 656.560 996.000 685.080 ;
        RECT 4.000 655.160 995.600 656.560 ;
        RECT 4.000 610.320 996.000 655.160 ;
        RECT 4.400 608.920 996.000 610.320 ;
        RECT 4.000 580.400 996.000 608.920 ;
        RECT 4.000 579.000 995.600 580.400 ;
        RECT 4.000 534.160 996.000 579.000 ;
        RECT 4.400 532.760 996.000 534.160 ;
        RECT 4.000 504.240 996.000 532.760 ;
        RECT 4.000 502.840 995.600 504.240 ;
        RECT 4.000 458.000 996.000 502.840 ;
        RECT 4.400 456.600 996.000 458.000 ;
        RECT 4.000 428.080 996.000 456.600 ;
        RECT 4.000 426.680 995.600 428.080 ;
        RECT 4.000 381.840 996.000 426.680 ;
        RECT 4.400 380.440 996.000 381.840 ;
        RECT 4.000 351.920 996.000 380.440 ;
        RECT 4.000 350.520 995.600 351.920 ;
        RECT 4.000 305.680 996.000 350.520 ;
        RECT 4.400 304.280 996.000 305.680 ;
        RECT 4.000 275.760 996.000 304.280 ;
        RECT 4.000 274.360 995.600 275.760 ;
        RECT 4.000 229.520 996.000 274.360 ;
        RECT 4.400 228.120 996.000 229.520 ;
        RECT 4.000 199.600 996.000 228.120 ;
        RECT 4.000 198.200 995.600 199.600 ;
        RECT 4.000 153.360 996.000 198.200 ;
        RECT 4.400 151.960 996.000 153.360 ;
        RECT 4.000 123.440 996.000 151.960 ;
        RECT 4.000 122.040 995.600 123.440 ;
        RECT 4.000 77.200 996.000 122.040 ;
        RECT 4.400 75.800 996.000 77.200 ;
        RECT 4.000 47.280 996.000 75.800 ;
        RECT 4.000 45.880 995.600 47.280 ;
        RECT 4.000 10.715 996.000 45.880 ;
  END
END multiplier
END LIBRARY

