magic
tech sky130A
magscale 1 2
timestamp 1641153771
<< metal1 >>
rect 211062 117988 211068 118040
rect 211120 118028 211126 118040
rect 284570 118028 284576 118040
rect 211120 118000 284576 118028
rect 211120 117988 211126 118000
rect 284570 117988 284576 118000
rect 284628 117988 284634 118040
rect 147582 117920 147588 117972
rect 147640 117960 147646 117972
rect 233234 117960 233240 117972
rect 147640 117932 233240 117960
rect 147640 117920 147646 117932
rect 233234 117920 233240 117932
rect 233292 117920 233298 117972
rect 151262 117308 151268 117360
rect 151320 117348 151326 117360
rect 151722 117348 151728 117360
rect 151320 117320 151728 117348
rect 151320 117308 151326 117320
rect 151722 117308 151728 117320
rect 151780 117308 151786 117360
rect 171870 117308 171876 117360
rect 171928 117348 171934 117360
rect 172422 117348 172428 117360
rect 171928 117320 172428 117348
rect 171928 117308 171934 117320
rect 172422 117308 172428 117320
rect 172480 117308 172486 117360
rect 118878 4088 118884 4140
rect 118936 4128 118942 4140
rect 164878 4128 164884 4140
rect 118936 4100 164884 4128
rect 118936 4088 118942 4100
rect 164878 4088 164884 4100
rect 164936 4088 164942 4140
rect 119982 4020 119988 4072
rect 120040 4060 120046 4072
rect 129366 4060 129372 4072
rect 120040 4032 129372 4060
rect 120040 4020 120046 4032
rect 129366 4020 129372 4032
rect 129424 4020 129430 4072
rect 140682 4020 140688 4072
rect 140740 4060 140746 4072
rect 193214 4060 193220 4072
rect 140740 4032 193220 4060
rect 140740 4020 140746 4032
rect 193214 4020 193220 4032
rect 193272 4020 193278 4072
rect 202782 4020 202788 4072
rect 202840 4060 202846 4072
rect 232222 4060 232228 4072
rect 202840 4032 232228 4060
rect 202840 4020 202846 4032
rect 232222 4020 232228 4032
rect 232280 4020 232286 4072
rect 118050 3952 118056 4004
rect 118108 3992 118114 4004
rect 171962 3992 171968 4004
rect 118108 3964 171968 3992
rect 118108 3952 118114 3964
rect 171962 3952 171968 3964
rect 172020 3952 172026 4004
rect 172422 3952 172428 4004
rect 172480 3992 172486 4004
rect 225138 3992 225144 4004
rect 172480 3964 225144 3992
rect 172480 3952 172486 3964
rect 225138 3952 225144 3964
rect 225196 3952 225202 4004
rect 118786 3884 118792 3936
rect 118844 3924 118850 3936
rect 132954 3924 132960 3936
rect 118844 3896 132960 3924
rect 118844 3884 118850 3896
rect 132954 3884 132960 3896
rect 133012 3884 133018 3936
rect 151722 3884 151728 3936
rect 151780 3924 151786 3936
rect 221550 3924 221556 3936
rect 151780 3896 221556 3924
rect 151780 3884 151786 3896
rect 221550 3884 221556 3896
rect 221608 3884 221614 3936
rect 118142 3816 118148 3868
rect 118200 3856 118206 3868
rect 214466 3856 214472 3868
rect 118200 3828 214472 3856
rect 118200 3816 118206 3828
rect 214466 3816 214472 3828
rect 214524 3816 214530 3868
rect 218054 3816 218060 3868
rect 218112 3856 218118 3868
rect 319070 3856 319076 3868
rect 218112 3828 319076 3856
rect 218112 3816 218118 3828
rect 319070 3816 319076 3828
rect 319128 3816 319134 3868
rect 118418 3748 118424 3800
rect 118476 3788 118482 3800
rect 228726 3788 228732 3800
rect 118476 3760 228732 3788
rect 118476 3748 118482 3760
rect 228726 3748 228732 3760
rect 228784 3748 228790 3800
rect 118510 3680 118516 3732
rect 118568 3720 118574 3732
rect 175458 3720 175464 3732
rect 118568 3692 175464 3720
rect 118568 3680 118574 3692
rect 175458 3680 175464 3692
rect 175516 3680 175522 3732
rect 182082 3680 182088 3732
rect 182140 3720 182146 3732
rect 203886 3720 203892 3732
rect 182140 3692 203892 3720
rect 182140 3680 182146 3692
rect 203886 3680 203892 3692
rect 203944 3680 203950 3732
rect 207382 3680 207388 3732
rect 207440 3720 207446 3732
rect 318886 3720 318892 3732
rect 207440 3692 318892 3720
rect 207440 3680 207446 3692
rect 318886 3680 318892 3692
rect 318944 3680 318950 3732
rect 118326 3612 118332 3664
rect 118384 3652 118390 3664
rect 182542 3652 182548 3664
rect 118384 3624 182548 3652
rect 118384 3612 118390 3624
rect 182542 3612 182548 3624
rect 182600 3612 182606 3664
rect 186130 3612 186136 3664
rect 186188 3652 186194 3664
rect 318794 3652 318800 3664
rect 186188 3624 318800 3652
rect 186188 3612 186194 3624
rect 318794 3612 318800 3624
rect 318852 3612 318858 3664
rect 118234 3544 118240 3596
rect 118292 3584 118298 3596
rect 150618 3584 150624 3596
rect 118292 3556 150624 3584
rect 118292 3544 118298 3556
rect 150618 3544 150624 3556
rect 150676 3544 150682 3596
rect 157794 3544 157800 3596
rect 157852 3584 157858 3596
rect 318978 3584 318984 3596
rect 157852 3556 318984 3584
rect 157852 3544 157858 3556
rect 318978 3544 318984 3556
rect 319036 3544 319042 3596
rect 125870 3476 125876 3528
rect 125928 3516 125934 3528
rect 319162 3516 319168 3528
rect 125928 3488 319168 3516
rect 125928 3476 125934 3488
rect 319162 3476 319168 3488
rect 319220 3476 319226 3528
rect 118602 3408 118608 3460
rect 118660 3448 118666 3460
rect 579798 3448 579804 3460
rect 118660 3420 579804 3448
rect 118660 3408 118666 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 147122 3340 147128 3392
rect 147180 3380 147186 3392
rect 147582 3380 147588 3392
rect 147180 3352 147588 3380
rect 147180 3340 147186 3352
rect 147582 3340 147588 3352
rect 147640 3340 147646 3392
<< via1 >>
rect 211068 117988 211120 118040
rect 284576 117988 284628 118040
rect 147588 117920 147640 117972
rect 233240 117920 233292 117972
rect 151268 117308 151320 117360
rect 151728 117308 151780 117360
rect 171876 117308 171928 117360
rect 172428 117308 172480 117360
rect 118884 4088 118936 4140
rect 164884 4088 164936 4140
rect 119988 4020 120040 4072
rect 129372 4020 129424 4072
rect 140688 4020 140740 4072
rect 193220 4020 193272 4072
rect 202788 4020 202840 4072
rect 232228 4020 232280 4072
rect 118056 3952 118108 4004
rect 171968 3952 172020 4004
rect 172428 3952 172480 4004
rect 225144 3952 225196 4004
rect 118792 3884 118844 3936
rect 132960 3884 133012 3936
rect 151728 3884 151780 3936
rect 221556 3884 221608 3936
rect 118148 3816 118200 3868
rect 214472 3816 214524 3868
rect 218060 3816 218112 3868
rect 319076 3816 319128 3868
rect 118424 3748 118476 3800
rect 228732 3748 228784 3800
rect 118516 3680 118568 3732
rect 175464 3680 175516 3732
rect 182088 3680 182140 3732
rect 203892 3680 203944 3732
rect 207388 3680 207440 3732
rect 318892 3680 318944 3732
rect 118332 3612 118384 3664
rect 182548 3612 182600 3664
rect 186136 3612 186188 3664
rect 318800 3612 318852 3664
rect 118240 3544 118292 3596
rect 150624 3544 150676 3596
rect 157800 3544 157852 3596
rect 318984 3544 319036 3596
rect 125876 3476 125928 3528
rect 319168 3476 319220 3528
rect 118608 3408 118660 3460
rect 579804 3408 579856 3460
rect 147128 3340 147180 3392
rect 147588 3340 147640 3392
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 139214 319424 139270 319433
rect 160466 319424 160522 319433
rect 139270 319382 139380 319410
rect 160172 319382 160466 319410
rect 139214 319359 139270 319368
rect 160466 319359 160522 319368
rect 170126 319424 170182 319433
rect 180430 319424 180486 319433
rect 170182 319382 170476 319410
rect 170126 319359 170182 319368
rect 201038 319424 201094 319433
rect 180486 319382 180780 319410
rect 180430 319359 180486 319368
rect 232594 319424 232650 319433
rect 201094 319382 201388 319410
rect 232300 319382 232594 319410
rect 201038 319359 201094 319368
rect 232594 319359 232650 319368
rect 273350 319424 273406 319433
rect 283470 319424 283526 319433
rect 273406 319382 273516 319410
rect 273350 319359 273406 319368
rect 293958 319424 294014 319433
rect 283526 319382 283820 319410
rect 283470 319359 283526 319368
rect 304078 319424 304134 319433
rect 294014 319382 294124 319410
rect 293958 319359 294014 319368
rect 314842 319424 314898 319433
rect 304134 319382 304428 319410
rect 314732 319382 314842 319410
rect 304078 319359 304134 319368
rect 314842 319359 314898 319368
rect 118514 287600 118570 287609
rect 118514 287535 118570 287544
rect 118422 257136 118478 257145
rect 118422 257071 118478 257080
rect 118330 241904 118386 241913
rect 118330 241839 118386 241848
rect 118238 211440 118294 211449
rect 118238 211375 118294 211384
rect 118146 196208 118202 196217
rect 118146 196143 118202 196152
rect 118054 150512 118110 150521
rect 118054 150447 118110 150456
rect 118068 4010 118096 150447
rect 118056 4004 118108 4010
rect 118056 3946 118108 3952
rect 118160 3874 118188 196143
rect 118148 3868 118200 3874
rect 118148 3810 118200 3816
rect 118252 3602 118280 211375
rect 118344 3670 118372 241839
rect 118436 3806 118464 257071
rect 118424 3800 118476 3806
rect 118424 3742 118476 3748
rect 118528 3738 118556 287535
rect 319350 281480 319406 281489
rect 319350 281415 319406 281424
rect 319364 277394 319392 281415
rect 318812 277366 319392 277394
rect 118606 272368 118662 272377
rect 118606 272303 118662 272312
rect 118516 3732 118568 3738
rect 118516 3674 118568 3680
rect 118332 3664 118384 3670
rect 118332 3606 118384 3612
rect 118240 3596 118292 3602
rect 118240 3538 118292 3544
rect 118620 3466 118648 272303
rect 118882 226672 118938 226681
rect 118882 226607 118938 226616
rect 118790 135280 118846 135289
rect 118790 135215 118846 135224
rect 118804 3942 118832 135215
rect 118896 4146 118924 226607
rect 120000 120006 120060 120034
rect 118884 4140 118936 4146
rect 118884 4082 118936 4088
rect 120000 4078 120028 120006
rect 140654 119762 140682 120020
rect 150972 120006 151308 120034
rect 171580 120006 171916 120034
rect 181884 120006 182128 120034
rect 202492 120006 202828 120034
rect 140654 119734 140728 119762
rect 140700 4078 140728 119734
rect 147588 117972 147640 117978
rect 147588 117914 147640 117920
rect 119988 4072 120040 4078
rect 119988 4014 120040 4020
rect 129372 4072 129424 4078
rect 129372 4014 129424 4020
rect 140688 4072 140740 4078
rect 140688 4014 140740 4020
rect 118792 3936 118844 3942
rect 118792 3878 118844 3884
rect 125876 3528 125928 3534
rect 125876 3470 125928 3476
rect 118608 3460 118660 3466
rect 118608 3402 118660 3408
rect 125888 480 125916 3470
rect 129384 480 129412 4014
rect 132960 3936 133012 3942
rect 132960 3878 133012 3884
rect 140042 3904 140098 3913
rect 132972 480 133000 3878
rect 140042 3839 140098 3848
rect 136454 3360 136510 3369
rect 136454 3295 136510 3304
rect 136468 480 136496 3295
rect 140056 480 140084 3839
rect 143538 3632 143594 3641
rect 143538 3567 143594 3576
rect 143552 480 143580 3567
rect 147600 3398 147628 117914
rect 151280 117366 151308 120006
rect 171888 117366 171916 120006
rect 151268 117360 151320 117366
rect 151268 117302 151320 117308
rect 151728 117360 151780 117366
rect 151728 117302 151780 117308
rect 171876 117360 171928 117366
rect 171876 117302 171928 117308
rect 172428 117360 172480 117366
rect 172428 117302 172480 117308
rect 151740 3942 151768 117302
rect 164884 4140 164936 4146
rect 164884 4082 164936 4088
rect 151728 3936 151780 3942
rect 151728 3878 151780 3884
rect 150624 3596 150676 3602
rect 150624 3538 150676 3544
rect 157800 3596 157852 3602
rect 157800 3538 157852 3544
rect 147128 3392 147180 3398
rect 147128 3334 147180 3340
rect 147588 3392 147640 3398
rect 147588 3334 147640 3340
rect 147140 480 147168 3334
rect 150636 480 150664 3538
rect 154210 3496 154266 3505
rect 154210 3431 154266 3440
rect 154224 480 154252 3431
rect 157812 480 157840 3538
rect 161294 3496 161350 3505
rect 161294 3431 161350 3440
rect 161308 480 161336 3431
rect 164896 480 164924 4082
rect 172440 4010 172468 117302
rect 171968 4004 172020 4010
rect 171968 3946 172020 3952
rect 172428 4004 172480 4010
rect 172428 3946 172480 3952
rect 168378 3768 168434 3777
rect 168378 3703 168434 3712
rect 168392 480 168420 3703
rect 171980 480 172008 3946
rect 179050 3768 179106 3777
rect 175464 3732 175516 3738
rect 182100 3738 182128 120006
rect 202800 4078 202828 120006
rect 233252 120006 233404 120034
rect 284588 120006 284924 120034
rect 211068 118040 211120 118046
rect 211068 117982 211120 117988
rect 211080 6914 211108 117982
rect 233252 117978 233280 120006
rect 284588 118046 284616 120006
rect 284576 118040 284628 118046
rect 284576 117982 284628 117988
rect 233240 117972 233292 117978
rect 233240 117914 233292 117920
rect 210988 6886 211108 6914
rect 193220 4072 193272 4078
rect 202788 4072 202840 4078
rect 193220 4014 193272 4020
rect 196806 4040 196862 4049
rect 189722 3904 189778 3913
rect 189722 3839 189778 3848
rect 179050 3703 179106 3712
rect 182088 3732 182140 3738
rect 175464 3674 175516 3680
rect 175476 480 175504 3674
rect 179064 480 179092 3703
rect 182088 3674 182140 3680
rect 182548 3664 182600 3670
rect 182548 3606 182600 3612
rect 186136 3664 186188 3670
rect 186136 3606 186188 3612
rect 182560 480 182588 3606
rect 186148 480 186176 3606
rect 189736 480 189764 3839
rect 193232 480 193260 4014
rect 202788 4014 202840 4020
rect 196806 3975 196862 3984
rect 196820 480 196848 3975
rect 203892 3732 203944 3738
rect 203892 3674 203944 3680
rect 207388 3732 207440 3738
rect 207388 3674 207440 3680
rect 200302 3632 200358 3641
rect 200302 3567 200358 3576
rect 200316 480 200344 3567
rect 203904 480 203932 3674
rect 207400 480 207428 3674
rect 210988 480 211016 6886
rect 232228 4072 232280 4078
rect 232228 4014 232280 4020
rect 225144 4004 225196 4010
rect 225144 3946 225196 3952
rect 221556 3936 221608 3942
rect 221556 3878 221608 3884
rect 214472 3868 214524 3874
rect 214472 3810 214524 3816
rect 218060 3868 218112 3874
rect 218060 3810 218112 3816
rect 214484 480 214512 3810
rect 218072 480 218100 3810
rect 221568 480 221596 3878
rect 225156 480 225184 3946
rect 228732 3800 228784 3806
rect 228732 3742 228784 3748
rect 228744 480 228772 3742
rect 232240 480 232268 4014
rect 235814 3904 235870 3913
rect 235814 3839 235870 3848
rect 235828 480 235856 3839
rect 318812 3670 318840 277366
rect 319350 266248 319406 266257
rect 319350 266183 319406 266192
rect 319364 258074 319392 266183
rect 318904 258046 319392 258074
rect 318904 3738 318932 258046
rect 319350 189680 319406 189689
rect 319350 189615 319406 189624
rect 319364 180794 319392 189615
rect 318996 180766 319392 180794
rect 318892 3732 318944 3738
rect 318892 3674 318944 3680
rect 318800 3664 318852 3670
rect 318800 3606 318852 3612
rect 318996 3602 319024 180766
rect 319350 174448 319406 174457
rect 319350 174383 319406 174392
rect 319364 161474 319392 174383
rect 319088 161446 319392 161474
rect 319088 3874 319116 161446
rect 319350 128752 319406 128761
rect 319350 128687 319406 128696
rect 319364 122834 319392 128687
rect 319180 122806 319392 122834
rect 319076 3868 319128 3874
rect 319076 3810 319128 3816
rect 318984 3596 319036 3602
rect 318984 3538 319036 3544
rect 319180 3534 319208 122806
rect 319168 3528 319220 3534
rect 319168 3470 319220 3476
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 139214 319368 139270 319424
rect 160466 319368 160522 319424
rect 170126 319368 170182 319424
rect 180430 319368 180486 319424
rect 201038 319368 201094 319424
rect 232594 319368 232650 319424
rect 273350 319368 273406 319424
rect 283470 319368 283526 319424
rect 293958 319368 294014 319424
rect 304078 319368 304134 319424
rect 314842 319368 314898 319424
rect 118514 287544 118570 287600
rect 118422 257080 118478 257136
rect 118330 241848 118386 241904
rect 118238 211384 118294 211440
rect 118146 196152 118202 196208
rect 118054 150456 118110 150512
rect 319350 281424 319406 281480
rect 118606 272312 118662 272368
rect 118882 226616 118938 226672
rect 118790 135224 118846 135280
rect 140042 3848 140098 3904
rect 136454 3304 136510 3360
rect 143538 3576 143594 3632
rect 154210 3440 154266 3496
rect 161294 3440 161350 3496
rect 168378 3712 168434 3768
rect 179050 3712 179106 3768
rect 189722 3848 189778 3904
rect 196806 3984 196862 4040
rect 200302 3576 200358 3632
rect 235814 3848 235870 3904
rect 319350 266192 319406 266248
rect 319350 189624 319406 189680
rect 319350 174392 319406 174448
rect 319350 128696 319406 128752
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect 139209 319428 139275 319429
rect 139158 319426 139164 319428
rect -960 319140 480 319380
rect 139118 319366 139164 319426
rect 139228 319424 139275 319428
rect 139270 319368 139275 319424
rect 139158 319364 139164 319366
rect 139228 319364 139275 319368
rect 139209 319363 139275 319364
rect 160461 319428 160527 319429
rect 160461 319424 160508 319428
rect 160572 319426 160578 319428
rect 160461 319368 160466 319424
rect 160461 319364 160508 319368
rect 160572 319366 160618 319426
rect 160572 319364 160578 319366
rect 169702 319364 169708 319428
rect 169772 319426 169778 319428
rect 170121 319426 170187 319429
rect 169772 319424 170187 319426
rect 169772 319368 170126 319424
rect 170182 319368 170187 319424
rect 169772 319366 170187 319368
rect 169772 319364 169778 319366
rect 160461 319363 160527 319364
rect 170121 319363 170187 319366
rect 179454 319364 179460 319428
rect 179524 319426 179530 319428
rect 180425 319426 180491 319429
rect 179524 319424 180491 319426
rect 179524 319368 180430 319424
rect 180486 319368 180491 319424
rect 179524 319366 180491 319368
rect 179524 319364 179530 319366
rect 180425 319363 180491 319366
rect 200246 319364 200252 319428
rect 200316 319426 200322 319428
rect 201033 319426 201099 319429
rect 200316 319424 201099 319426
rect 200316 319368 201038 319424
rect 201094 319368 201099 319424
rect 200316 319366 201099 319368
rect 200316 319364 200322 319366
rect 201033 319363 201099 319366
rect 232589 319426 232655 319429
rect 273345 319428 273411 319429
rect 232814 319426 232820 319428
rect 232589 319424 232820 319426
rect 232589 319368 232594 319424
rect 232650 319368 232820 319424
rect 232589 319366 232820 319368
rect 232589 319363 232655 319366
rect 232814 319364 232820 319366
rect 232884 319364 232890 319428
rect 273294 319426 273300 319428
rect 273254 319366 273300 319426
rect 273364 319424 273411 319428
rect 273406 319368 273411 319424
rect 273294 319364 273300 319366
rect 273364 319364 273411 319368
rect 282862 319364 282868 319428
rect 282932 319426 282938 319428
rect 283465 319426 283531 319429
rect 293953 319428 294019 319429
rect 293902 319426 293908 319428
rect 282932 319424 283531 319426
rect 282932 319368 283470 319424
rect 283526 319368 283531 319424
rect 282932 319366 283531 319368
rect 293862 319366 293908 319426
rect 293972 319424 294019 319428
rect 294014 319368 294019 319424
rect 282932 319364 282938 319366
rect 273345 319363 273411 319364
rect 283465 319363 283531 319366
rect 293902 319364 293908 319366
rect 293972 319364 294019 319368
rect 303654 319364 303660 319428
rect 303724 319426 303730 319428
rect 304073 319426 304139 319429
rect 303724 319424 304139 319426
rect 303724 319368 304078 319424
rect 304134 319368 304139 319424
rect 303724 319366 304139 319368
rect 303724 319364 303730 319366
rect 293953 319363 294019 319364
rect 304073 319363 304139 319366
rect 314694 319364 314700 319428
rect 314764 319426 314770 319428
rect 314837 319426 314903 319429
rect 314764 319424 314903 319426
rect 314764 319368 314842 319424
rect 314898 319368 314903 319424
rect 314764 319366 314903 319368
rect 314764 319364 314770 319366
rect 314837 319363 314903 319366
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 118509 287602 118575 287605
rect 118509 287600 120060 287602
rect 118509 287544 118514 287600
rect 118570 287544 120060 287600
rect 118509 287542 120060 287544
rect 118509 287539 118575 287542
rect 583520 285276 584960 285516
rect 319302 281485 319362 281588
rect 319302 281480 319411 281485
rect 319302 281424 319350 281480
rect 319406 281424 319411 281480
rect 319302 281422 319411 281424
rect 319345 281419 319411 281422
rect -960 279972 480 280212
rect 118601 272370 118667 272373
rect 118601 272368 120060 272370
rect 118601 272312 118606 272368
rect 118662 272312 120060 272368
rect 118601 272310 120060 272312
rect 118601 272307 118667 272310
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 319302 266253 319362 266356
rect 319302 266248 319411 266253
rect 319302 266192 319350 266248
rect 319406 266192 319411 266248
rect 319302 266190 319411 266192
rect 319345 266187 319411 266190
rect 583520 258756 584960 258996
rect 118417 257138 118483 257141
rect 118417 257136 120060 257138
rect 118417 257080 118422 257136
rect 118478 257080 120060 257136
rect 118417 257078 120060 257080
rect 118417 257075 118483 257078
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect 118325 241906 118391 241909
rect 118325 241904 120060 241906
rect 118325 241848 118330 241904
rect 118386 241848 120060 241904
rect 118325 241846 120060 241848
rect 118325 241843 118391 241846
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 118877 226674 118943 226677
rect 118877 226672 120060 226674
rect 118877 226616 118882 226672
rect 118938 226616 120060 226672
rect 118877 226614 120060 226616
rect 118877 226611 118943 226614
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 118233 211442 118299 211445
rect 118233 211440 120060 211442
rect 118233 211384 118238 211440
rect 118294 211384 120060 211440
rect 118233 211382 120060 211384
rect 118233 211379 118299 211382
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 118141 196210 118207 196213
rect 118141 196208 120060 196210
rect 118141 196152 118146 196208
rect 118202 196152 120060 196208
rect 118141 196150 120060 196152
rect 118141 196147 118207 196150
rect 583520 192388 584960 192628
rect 319302 189685 319362 190196
rect 319302 189680 319411 189685
rect 319302 189624 319350 189680
rect 319406 189624 319411 189680
rect 319302 189622 319411 189624
rect 319345 189619 319411 189622
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 319302 174453 319362 174964
rect 319302 174448 319411 174453
rect 319302 174392 319350 174448
rect 319406 174392 319411 174448
rect 319302 174390 319411 174392
rect 319345 174387 319411 174390
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect 118049 150514 118115 150517
rect 118049 150512 120060 150514
rect 118049 150456 118054 150512
rect 118110 150456 120060 150512
rect 118049 150454 120060 150456
rect 118049 150451 118115 150454
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 118785 135282 118851 135285
rect 118785 135280 120060 135282
rect 118785 135224 118790 135280
rect 118846 135224 120060 135280
rect 118785 135222 120060 135224
rect 118785 135219 118851 135222
rect 319302 128757 319362 129268
rect 319302 128752 319411 128757
rect 319302 128696 319350 128752
rect 319406 128696 319411 128752
rect 319302 128694 319411 128696
rect 319345 128691 319411 128694
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 160502 3980 160508 4044
rect 160572 4042 160578 4044
rect 196801 4042 196867 4045
rect 160572 4040 196867 4042
rect 160572 3984 196806 4040
rect 196862 3984 196867 4040
rect 160572 3982 196867 3984
rect 160572 3980 160578 3982
rect 196801 3979 196867 3982
rect 140037 3906 140103 3909
rect 179454 3906 179460 3908
rect 140037 3904 179460 3906
rect 140037 3848 140042 3904
rect 140098 3848 179460 3904
rect 140037 3846 179460 3848
rect 140037 3843 140103 3846
rect 179454 3844 179460 3846
rect 179524 3844 179530 3908
rect 189717 3906 189783 3909
rect 232814 3906 232820 3908
rect 189717 3904 232820 3906
rect 189717 3848 189722 3904
rect 189778 3848 232820 3904
rect 189717 3846 232820 3848
rect 189717 3843 189783 3846
rect 232814 3844 232820 3846
rect 232884 3844 232890 3908
rect 235809 3906 235875 3909
rect 303654 3906 303660 3908
rect 235809 3904 303660 3906
rect 235809 3848 235814 3904
rect 235870 3848 303660 3904
rect 235809 3846 303660 3848
rect 235809 3843 235875 3846
rect 303654 3844 303660 3846
rect 303724 3844 303730 3908
rect 168373 3770 168439 3773
rect 169702 3770 169708 3772
rect 168373 3768 169708 3770
rect 168373 3712 168378 3768
rect 168434 3712 169708 3768
rect 168373 3710 169708 3712
rect 168373 3707 168439 3710
rect 169702 3708 169708 3710
rect 169772 3708 169778 3772
rect 179045 3770 179111 3773
rect 273294 3770 273300 3772
rect 179045 3768 273300 3770
rect 179045 3712 179050 3768
rect 179106 3712 273300 3768
rect 179045 3710 273300 3712
rect 179045 3707 179111 3710
rect 273294 3708 273300 3710
rect 273364 3708 273370 3772
rect 143533 3634 143599 3637
rect 199878 3634 199884 3636
rect 143533 3632 199884 3634
rect 143533 3576 143538 3632
rect 143594 3576 199884 3632
rect 143533 3574 199884 3576
rect 143533 3571 143599 3574
rect 199878 3572 199884 3574
rect 199948 3572 199954 3636
rect 200297 3634 200363 3637
rect 314694 3634 314700 3636
rect 200297 3632 314700 3634
rect 200297 3576 200302 3632
rect 200358 3576 314700 3632
rect 200297 3574 314700 3576
rect 200297 3571 200363 3574
rect 314694 3572 314700 3574
rect 314764 3572 314770 3636
rect 139158 3436 139164 3500
rect 139228 3498 139234 3500
rect 154205 3498 154271 3501
rect 139228 3496 154271 3498
rect 139228 3440 154210 3496
rect 154266 3440 154271 3496
rect 139228 3438 154271 3440
rect 139228 3436 139234 3438
rect 154205 3435 154271 3438
rect 161289 3498 161355 3501
rect 282862 3498 282868 3500
rect 161289 3496 282868 3498
rect 161289 3440 161294 3496
rect 161350 3440 282868 3496
rect 161289 3438 282868 3440
rect 161289 3435 161355 3438
rect 282862 3436 282868 3438
rect 282932 3436 282938 3500
rect 136449 3362 136515 3365
rect 293902 3362 293908 3364
rect 136449 3360 293908 3362
rect 136449 3304 136454 3360
rect 136510 3304 293908 3360
rect 136449 3302 293908 3304
rect 136449 3299 136515 3302
rect 293902 3300 293908 3302
rect 293972 3300 293978 3364
<< via3 >>
rect 139164 319424 139228 319428
rect 139164 319368 139214 319424
rect 139214 319368 139228 319424
rect 139164 319364 139228 319368
rect 160508 319424 160572 319428
rect 160508 319368 160522 319424
rect 160522 319368 160572 319424
rect 160508 319364 160572 319368
rect 169708 319364 169772 319428
rect 179460 319364 179524 319428
rect 200252 319364 200316 319428
rect 232820 319364 232884 319428
rect 273300 319424 273364 319428
rect 273300 319368 273350 319424
rect 273350 319368 273364 319424
rect 273300 319364 273364 319368
rect 282868 319364 282932 319428
rect 293908 319424 293972 319428
rect 293908 319368 293958 319424
rect 293958 319368 293972 319424
rect 293908 319364 293972 319368
rect 303660 319364 303724 319428
rect 314700 319364 314764 319428
rect 160508 3980 160572 4044
rect 179460 3844 179524 3908
rect 232820 3844 232884 3908
rect 303660 3844 303724 3908
rect 169708 3708 169772 3772
rect 273300 3708 273364 3772
rect 199884 3572 199948 3636
rect 314700 3572 314764 3636
rect 139164 3436 139228 3500
rect 282868 3436 282932 3500
rect 293908 3300 293972 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 673614 -8106 711002
rect -8726 673378 -8694 673614
rect -8458 673378 -8374 673614
rect -8138 673378 -8106 673614
rect -8726 673294 -8106 673378
rect -8726 673058 -8694 673294
rect -8458 673058 -8374 673294
rect -8138 673058 -8106 673294
rect -8726 633614 -8106 673058
rect -8726 633378 -8694 633614
rect -8458 633378 -8374 633614
rect -8138 633378 -8106 633614
rect -8726 633294 -8106 633378
rect -8726 633058 -8694 633294
rect -8458 633058 -8374 633294
rect -8138 633058 -8106 633294
rect -8726 593614 -8106 633058
rect -8726 593378 -8694 593614
rect -8458 593378 -8374 593614
rect -8138 593378 -8106 593614
rect -8726 593294 -8106 593378
rect -8726 593058 -8694 593294
rect -8458 593058 -8374 593294
rect -8138 593058 -8106 593294
rect -8726 553614 -8106 593058
rect -8726 553378 -8694 553614
rect -8458 553378 -8374 553614
rect -8138 553378 -8106 553614
rect -8726 553294 -8106 553378
rect -8726 553058 -8694 553294
rect -8458 553058 -8374 553294
rect -8138 553058 -8106 553294
rect -8726 513614 -8106 553058
rect -8726 513378 -8694 513614
rect -8458 513378 -8374 513614
rect -8138 513378 -8106 513614
rect -8726 513294 -8106 513378
rect -8726 513058 -8694 513294
rect -8458 513058 -8374 513294
rect -8138 513058 -8106 513294
rect -8726 473614 -8106 513058
rect -8726 473378 -8694 473614
rect -8458 473378 -8374 473614
rect -8138 473378 -8106 473614
rect -8726 473294 -8106 473378
rect -8726 473058 -8694 473294
rect -8458 473058 -8374 473294
rect -8138 473058 -8106 473294
rect -8726 433614 -8106 473058
rect -8726 433378 -8694 433614
rect -8458 433378 -8374 433614
rect -8138 433378 -8106 433614
rect -8726 433294 -8106 433378
rect -8726 433058 -8694 433294
rect -8458 433058 -8374 433294
rect -8138 433058 -8106 433294
rect -8726 393614 -8106 433058
rect -8726 393378 -8694 393614
rect -8458 393378 -8374 393614
rect -8138 393378 -8106 393614
rect -8726 393294 -8106 393378
rect -8726 393058 -8694 393294
rect -8458 393058 -8374 393294
rect -8138 393058 -8106 393294
rect -8726 353614 -8106 393058
rect -8726 353378 -8694 353614
rect -8458 353378 -8374 353614
rect -8138 353378 -8106 353614
rect -8726 353294 -8106 353378
rect -8726 353058 -8694 353294
rect -8458 353058 -8374 353294
rect -8138 353058 -8106 353294
rect -8726 313614 -8106 353058
rect -8726 313378 -8694 313614
rect -8458 313378 -8374 313614
rect -8138 313378 -8106 313614
rect -8726 313294 -8106 313378
rect -8726 313058 -8694 313294
rect -8458 313058 -8374 313294
rect -8138 313058 -8106 313294
rect -8726 273614 -8106 313058
rect -8726 273378 -8694 273614
rect -8458 273378 -8374 273614
rect -8138 273378 -8106 273614
rect -8726 273294 -8106 273378
rect -8726 273058 -8694 273294
rect -8458 273058 -8374 273294
rect -8138 273058 -8106 273294
rect -8726 233614 -8106 273058
rect -8726 233378 -8694 233614
rect -8458 233378 -8374 233614
rect -8138 233378 -8106 233614
rect -8726 233294 -8106 233378
rect -8726 233058 -8694 233294
rect -8458 233058 -8374 233294
rect -8138 233058 -8106 233294
rect -8726 193614 -8106 233058
rect -8726 193378 -8694 193614
rect -8458 193378 -8374 193614
rect -8138 193378 -8106 193614
rect -8726 193294 -8106 193378
rect -8726 193058 -8694 193294
rect -8458 193058 -8374 193294
rect -8138 193058 -8106 193294
rect -8726 153614 -8106 193058
rect -8726 153378 -8694 153614
rect -8458 153378 -8374 153614
rect -8138 153378 -8106 153614
rect -8726 153294 -8106 153378
rect -8726 153058 -8694 153294
rect -8458 153058 -8374 153294
rect -8138 153058 -8106 153294
rect -8726 113614 -8106 153058
rect -8726 113378 -8694 113614
rect -8458 113378 -8374 113614
rect -8138 113378 -8106 113614
rect -8726 113294 -8106 113378
rect -8726 113058 -8694 113294
rect -8458 113058 -8374 113294
rect -8138 113058 -8106 113294
rect -8726 73614 -8106 113058
rect -8726 73378 -8694 73614
rect -8458 73378 -8374 73614
rect -8138 73378 -8106 73614
rect -8726 73294 -8106 73378
rect -8726 73058 -8694 73294
rect -8458 73058 -8374 73294
rect -8138 73058 -8106 73294
rect -8726 33614 -8106 73058
rect -8726 33378 -8694 33614
rect -8458 33378 -8374 33614
rect -8138 33378 -8106 33614
rect -8726 33294 -8106 33378
rect -8726 33058 -8694 33294
rect -8458 33058 -8374 33294
rect -8138 33058 -8106 33294
rect -8726 -7066 -8106 33058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 693614 -7146 710042
rect 11954 710598 12574 711590
rect 11954 710362 11986 710598
rect 12222 710362 12306 710598
rect 12542 710362 12574 710598
rect 11954 710278 12574 710362
rect 11954 710042 11986 710278
rect 12222 710042 12306 710278
rect 12542 710042 12574 710278
rect -7766 693378 -7734 693614
rect -7498 693378 -7414 693614
rect -7178 693378 -7146 693614
rect -7766 693294 -7146 693378
rect -7766 693058 -7734 693294
rect -7498 693058 -7414 693294
rect -7178 693058 -7146 693294
rect -7766 653614 -7146 693058
rect -7766 653378 -7734 653614
rect -7498 653378 -7414 653614
rect -7178 653378 -7146 653614
rect -7766 653294 -7146 653378
rect -7766 653058 -7734 653294
rect -7498 653058 -7414 653294
rect -7178 653058 -7146 653294
rect -7766 613614 -7146 653058
rect -7766 613378 -7734 613614
rect -7498 613378 -7414 613614
rect -7178 613378 -7146 613614
rect -7766 613294 -7146 613378
rect -7766 613058 -7734 613294
rect -7498 613058 -7414 613294
rect -7178 613058 -7146 613294
rect -7766 573614 -7146 613058
rect -7766 573378 -7734 573614
rect -7498 573378 -7414 573614
rect -7178 573378 -7146 573614
rect -7766 573294 -7146 573378
rect -7766 573058 -7734 573294
rect -7498 573058 -7414 573294
rect -7178 573058 -7146 573294
rect -7766 533614 -7146 573058
rect -7766 533378 -7734 533614
rect -7498 533378 -7414 533614
rect -7178 533378 -7146 533614
rect -7766 533294 -7146 533378
rect -7766 533058 -7734 533294
rect -7498 533058 -7414 533294
rect -7178 533058 -7146 533294
rect -7766 493614 -7146 533058
rect -7766 493378 -7734 493614
rect -7498 493378 -7414 493614
rect -7178 493378 -7146 493614
rect -7766 493294 -7146 493378
rect -7766 493058 -7734 493294
rect -7498 493058 -7414 493294
rect -7178 493058 -7146 493294
rect -7766 453614 -7146 493058
rect -7766 453378 -7734 453614
rect -7498 453378 -7414 453614
rect -7178 453378 -7146 453614
rect -7766 453294 -7146 453378
rect -7766 453058 -7734 453294
rect -7498 453058 -7414 453294
rect -7178 453058 -7146 453294
rect -7766 413614 -7146 453058
rect -7766 413378 -7734 413614
rect -7498 413378 -7414 413614
rect -7178 413378 -7146 413614
rect -7766 413294 -7146 413378
rect -7766 413058 -7734 413294
rect -7498 413058 -7414 413294
rect -7178 413058 -7146 413294
rect -7766 373614 -7146 413058
rect -7766 373378 -7734 373614
rect -7498 373378 -7414 373614
rect -7178 373378 -7146 373614
rect -7766 373294 -7146 373378
rect -7766 373058 -7734 373294
rect -7498 373058 -7414 373294
rect -7178 373058 -7146 373294
rect -7766 333614 -7146 373058
rect -7766 333378 -7734 333614
rect -7498 333378 -7414 333614
rect -7178 333378 -7146 333614
rect -7766 333294 -7146 333378
rect -7766 333058 -7734 333294
rect -7498 333058 -7414 333294
rect -7178 333058 -7146 333294
rect -7766 293614 -7146 333058
rect -7766 293378 -7734 293614
rect -7498 293378 -7414 293614
rect -7178 293378 -7146 293614
rect -7766 293294 -7146 293378
rect -7766 293058 -7734 293294
rect -7498 293058 -7414 293294
rect -7178 293058 -7146 293294
rect -7766 253614 -7146 293058
rect -7766 253378 -7734 253614
rect -7498 253378 -7414 253614
rect -7178 253378 -7146 253614
rect -7766 253294 -7146 253378
rect -7766 253058 -7734 253294
rect -7498 253058 -7414 253294
rect -7178 253058 -7146 253294
rect -7766 213614 -7146 253058
rect -7766 213378 -7734 213614
rect -7498 213378 -7414 213614
rect -7178 213378 -7146 213614
rect -7766 213294 -7146 213378
rect -7766 213058 -7734 213294
rect -7498 213058 -7414 213294
rect -7178 213058 -7146 213294
rect -7766 173614 -7146 213058
rect -7766 173378 -7734 173614
rect -7498 173378 -7414 173614
rect -7178 173378 -7146 173614
rect -7766 173294 -7146 173378
rect -7766 173058 -7734 173294
rect -7498 173058 -7414 173294
rect -7178 173058 -7146 173294
rect -7766 133614 -7146 173058
rect -7766 133378 -7734 133614
rect -7498 133378 -7414 133614
rect -7178 133378 -7146 133614
rect -7766 133294 -7146 133378
rect -7766 133058 -7734 133294
rect -7498 133058 -7414 133294
rect -7178 133058 -7146 133294
rect -7766 93614 -7146 133058
rect -7766 93378 -7734 93614
rect -7498 93378 -7414 93614
rect -7178 93378 -7146 93614
rect -7766 93294 -7146 93378
rect -7766 93058 -7734 93294
rect -7498 93058 -7414 93294
rect -7178 93058 -7146 93294
rect -7766 53614 -7146 93058
rect -7766 53378 -7734 53614
rect -7498 53378 -7414 53614
rect -7178 53378 -7146 53614
rect -7766 53294 -7146 53378
rect -7766 53058 -7734 53294
rect -7498 53058 -7414 53294
rect -7178 53058 -7146 53294
rect -7766 13614 -7146 53058
rect -7766 13378 -7734 13614
rect -7498 13378 -7414 13614
rect -7178 13378 -7146 13614
rect -7766 13294 -7146 13378
rect -7766 13058 -7734 13294
rect -7498 13058 -7414 13294
rect -7178 13058 -7146 13294
rect -7766 -6106 -7146 13058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 669894 -6186 709082
rect -6806 669658 -6774 669894
rect -6538 669658 -6454 669894
rect -6218 669658 -6186 669894
rect -6806 669574 -6186 669658
rect -6806 669338 -6774 669574
rect -6538 669338 -6454 669574
rect -6218 669338 -6186 669574
rect -6806 629894 -6186 669338
rect -6806 629658 -6774 629894
rect -6538 629658 -6454 629894
rect -6218 629658 -6186 629894
rect -6806 629574 -6186 629658
rect -6806 629338 -6774 629574
rect -6538 629338 -6454 629574
rect -6218 629338 -6186 629574
rect -6806 589894 -6186 629338
rect -6806 589658 -6774 589894
rect -6538 589658 -6454 589894
rect -6218 589658 -6186 589894
rect -6806 589574 -6186 589658
rect -6806 589338 -6774 589574
rect -6538 589338 -6454 589574
rect -6218 589338 -6186 589574
rect -6806 549894 -6186 589338
rect -6806 549658 -6774 549894
rect -6538 549658 -6454 549894
rect -6218 549658 -6186 549894
rect -6806 549574 -6186 549658
rect -6806 549338 -6774 549574
rect -6538 549338 -6454 549574
rect -6218 549338 -6186 549574
rect -6806 509894 -6186 549338
rect -6806 509658 -6774 509894
rect -6538 509658 -6454 509894
rect -6218 509658 -6186 509894
rect -6806 509574 -6186 509658
rect -6806 509338 -6774 509574
rect -6538 509338 -6454 509574
rect -6218 509338 -6186 509574
rect -6806 469894 -6186 509338
rect -6806 469658 -6774 469894
rect -6538 469658 -6454 469894
rect -6218 469658 -6186 469894
rect -6806 469574 -6186 469658
rect -6806 469338 -6774 469574
rect -6538 469338 -6454 469574
rect -6218 469338 -6186 469574
rect -6806 429894 -6186 469338
rect -6806 429658 -6774 429894
rect -6538 429658 -6454 429894
rect -6218 429658 -6186 429894
rect -6806 429574 -6186 429658
rect -6806 429338 -6774 429574
rect -6538 429338 -6454 429574
rect -6218 429338 -6186 429574
rect -6806 389894 -6186 429338
rect -6806 389658 -6774 389894
rect -6538 389658 -6454 389894
rect -6218 389658 -6186 389894
rect -6806 389574 -6186 389658
rect -6806 389338 -6774 389574
rect -6538 389338 -6454 389574
rect -6218 389338 -6186 389574
rect -6806 349894 -6186 389338
rect -6806 349658 -6774 349894
rect -6538 349658 -6454 349894
rect -6218 349658 -6186 349894
rect -6806 349574 -6186 349658
rect -6806 349338 -6774 349574
rect -6538 349338 -6454 349574
rect -6218 349338 -6186 349574
rect -6806 309894 -6186 349338
rect -6806 309658 -6774 309894
rect -6538 309658 -6454 309894
rect -6218 309658 -6186 309894
rect -6806 309574 -6186 309658
rect -6806 309338 -6774 309574
rect -6538 309338 -6454 309574
rect -6218 309338 -6186 309574
rect -6806 269894 -6186 309338
rect -6806 269658 -6774 269894
rect -6538 269658 -6454 269894
rect -6218 269658 -6186 269894
rect -6806 269574 -6186 269658
rect -6806 269338 -6774 269574
rect -6538 269338 -6454 269574
rect -6218 269338 -6186 269574
rect -6806 229894 -6186 269338
rect -6806 229658 -6774 229894
rect -6538 229658 -6454 229894
rect -6218 229658 -6186 229894
rect -6806 229574 -6186 229658
rect -6806 229338 -6774 229574
rect -6538 229338 -6454 229574
rect -6218 229338 -6186 229574
rect -6806 189894 -6186 229338
rect -6806 189658 -6774 189894
rect -6538 189658 -6454 189894
rect -6218 189658 -6186 189894
rect -6806 189574 -6186 189658
rect -6806 189338 -6774 189574
rect -6538 189338 -6454 189574
rect -6218 189338 -6186 189574
rect -6806 149894 -6186 189338
rect -6806 149658 -6774 149894
rect -6538 149658 -6454 149894
rect -6218 149658 -6186 149894
rect -6806 149574 -6186 149658
rect -6806 149338 -6774 149574
rect -6538 149338 -6454 149574
rect -6218 149338 -6186 149574
rect -6806 109894 -6186 149338
rect -6806 109658 -6774 109894
rect -6538 109658 -6454 109894
rect -6218 109658 -6186 109894
rect -6806 109574 -6186 109658
rect -6806 109338 -6774 109574
rect -6538 109338 -6454 109574
rect -6218 109338 -6186 109574
rect -6806 69894 -6186 109338
rect -6806 69658 -6774 69894
rect -6538 69658 -6454 69894
rect -6218 69658 -6186 69894
rect -6806 69574 -6186 69658
rect -6806 69338 -6774 69574
rect -6538 69338 -6454 69574
rect -6218 69338 -6186 69574
rect -6806 29894 -6186 69338
rect -6806 29658 -6774 29894
rect -6538 29658 -6454 29894
rect -6218 29658 -6186 29894
rect -6806 29574 -6186 29658
rect -6806 29338 -6774 29574
rect -6538 29338 -6454 29574
rect -6218 29338 -6186 29574
rect -6806 -5146 -6186 29338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 689894 -5226 708122
rect 8234 708678 8854 709670
rect 8234 708442 8266 708678
rect 8502 708442 8586 708678
rect 8822 708442 8854 708678
rect 8234 708358 8854 708442
rect 8234 708122 8266 708358
rect 8502 708122 8586 708358
rect 8822 708122 8854 708358
rect -5846 689658 -5814 689894
rect -5578 689658 -5494 689894
rect -5258 689658 -5226 689894
rect -5846 689574 -5226 689658
rect -5846 689338 -5814 689574
rect -5578 689338 -5494 689574
rect -5258 689338 -5226 689574
rect -5846 649894 -5226 689338
rect -5846 649658 -5814 649894
rect -5578 649658 -5494 649894
rect -5258 649658 -5226 649894
rect -5846 649574 -5226 649658
rect -5846 649338 -5814 649574
rect -5578 649338 -5494 649574
rect -5258 649338 -5226 649574
rect -5846 609894 -5226 649338
rect -5846 609658 -5814 609894
rect -5578 609658 -5494 609894
rect -5258 609658 -5226 609894
rect -5846 609574 -5226 609658
rect -5846 609338 -5814 609574
rect -5578 609338 -5494 609574
rect -5258 609338 -5226 609574
rect -5846 569894 -5226 609338
rect -5846 569658 -5814 569894
rect -5578 569658 -5494 569894
rect -5258 569658 -5226 569894
rect -5846 569574 -5226 569658
rect -5846 569338 -5814 569574
rect -5578 569338 -5494 569574
rect -5258 569338 -5226 569574
rect -5846 529894 -5226 569338
rect -5846 529658 -5814 529894
rect -5578 529658 -5494 529894
rect -5258 529658 -5226 529894
rect -5846 529574 -5226 529658
rect -5846 529338 -5814 529574
rect -5578 529338 -5494 529574
rect -5258 529338 -5226 529574
rect -5846 489894 -5226 529338
rect -5846 489658 -5814 489894
rect -5578 489658 -5494 489894
rect -5258 489658 -5226 489894
rect -5846 489574 -5226 489658
rect -5846 489338 -5814 489574
rect -5578 489338 -5494 489574
rect -5258 489338 -5226 489574
rect -5846 449894 -5226 489338
rect -5846 449658 -5814 449894
rect -5578 449658 -5494 449894
rect -5258 449658 -5226 449894
rect -5846 449574 -5226 449658
rect -5846 449338 -5814 449574
rect -5578 449338 -5494 449574
rect -5258 449338 -5226 449574
rect -5846 409894 -5226 449338
rect -5846 409658 -5814 409894
rect -5578 409658 -5494 409894
rect -5258 409658 -5226 409894
rect -5846 409574 -5226 409658
rect -5846 409338 -5814 409574
rect -5578 409338 -5494 409574
rect -5258 409338 -5226 409574
rect -5846 369894 -5226 409338
rect -5846 369658 -5814 369894
rect -5578 369658 -5494 369894
rect -5258 369658 -5226 369894
rect -5846 369574 -5226 369658
rect -5846 369338 -5814 369574
rect -5578 369338 -5494 369574
rect -5258 369338 -5226 369574
rect -5846 329894 -5226 369338
rect -5846 329658 -5814 329894
rect -5578 329658 -5494 329894
rect -5258 329658 -5226 329894
rect -5846 329574 -5226 329658
rect -5846 329338 -5814 329574
rect -5578 329338 -5494 329574
rect -5258 329338 -5226 329574
rect -5846 289894 -5226 329338
rect -5846 289658 -5814 289894
rect -5578 289658 -5494 289894
rect -5258 289658 -5226 289894
rect -5846 289574 -5226 289658
rect -5846 289338 -5814 289574
rect -5578 289338 -5494 289574
rect -5258 289338 -5226 289574
rect -5846 249894 -5226 289338
rect -5846 249658 -5814 249894
rect -5578 249658 -5494 249894
rect -5258 249658 -5226 249894
rect -5846 249574 -5226 249658
rect -5846 249338 -5814 249574
rect -5578 249338 -5494 249574
rect -5258 249338 -5226 249574
rect -5846 209894 -5226 249338
rect -5846 209658 -5814 209894
rect -5578 209658 -5494 209894
rect -5258 209658 -5226 209894
rect -5846 209574 -5226 209658
rect -5846 209338 -5814 209574
rect -5578 209338 -5494 209574
rect -5258 209338 -5226 209574
rect -5846 169894 -5226 209338
rect -5846 169658 -5814 169894
rect -5578 169658 -5494 169894
rect -5258 169658 -5226 169894
rect -5846 169574 -5226 169658
rect -5846 169338 -5814 169574
rect -5578 169338 -5494 169574
rect -5258 169338 -5226 169574
rect -5846 129894 -5226 169338
rect -5846 129658 -5814 129894
rect -5578 129658 -5494 129894
rect -5258 129658 -5226 129894
rect -5846 129574 -5226 129658
rect -5846 129338 -5814 129574
rect -5578 129338 -5494 129574
rect -5258 129338 -5226 129574
rect -5846 89894 -5226 129338
rect -5846 89658 -5814 89894
rect -5578 89658 -5494 89894
rect -5258 89658 -5226 89894
rect -5846 89574 -5226 89658
rect -5846 89338 -5814 89574
rect -5578 89338 -5494 89574
rect -5258 89338 -5226 89574
rect -5846 49894 -5226 89338
rect -5846 49658 -5814 49894
rect -5578 49658 -5494 49894
rect -5258 49658 -5226 49894
rect -5846 49574 -5226 49658
rect -5846 49338 -5814 49574
rect -5578 49338 -5494 49574
rect -5258 49338 -5226 49574
rect -5846 9894 -5226 49338
rect -5846 9658 -5814 9894
rect -5578 9658 -5494 9894
rect -5258 9658 -5226 9894
rect -5846 9574 -5226 9658
rect -5846 9338 -5814 9574
rect -5578 9338 -5494 9574
rect -5258 9338 -5226 9574
rect -5846 -4186 -5226 9338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 666174 -4266 707162
rect -4886 665938 -4854 666174
rect -4618 665938 -4534 666174
rect -4298 665938 -4266 666174
rect -4886 665854 -4266 665938
rect -4886 665618 -4854 665854
rect -4618 665618 -4534 665854
rect -4298 665618 -4266 665854
rect -4886 626174 -4266 665618
rect -4886 625938 -4854 626174
rect -4618 625938 -4534 626174
rect -4298 625938 -4266 626174
rect -4886 625854 -4266 625938
rect -4886 625618 -4854 625854
rect -4618 625618 -4534 625854
rect -4298 625618 -4266 625854
rect -4886 586174 -4266 625618
rect -4886 585938 -4854 586174
rect -4618 585938 -4534 586174
rect -4298 585938 -4266 586174
rect -4886 585854 -4266 585938
rect -4886 585618 -4854 585854
rect -4618 585618 -4534 585854
rect -4298 585618 -4266 585854
rect -4886 546174 -4266 585618
rect -4886 545938 -4854 546174
rect -4618 545938 -4534 546174
rect -4298 545938 -4266 546174
rect -4886 545854 -4266 545938
rect -4886 545618 -4854 545854
rect -4618 545618 -4534 545854
rect -4298 545618 -4266 545854
rect -4886 506174 -4266 545618
rect -4886 505938 -4854 506174
rect -4618 505938 -4534 506174
rect -4298 505938 -4266 506174
rect -4886 505854 -4266 505938
rect -4886 505618 -4854 505854
rect -4618 505618 -4534 505854
rect -4298 505618 -4266 505854
rect -4886 466174 -4266 505618
rect -4886 465938 -4854 466174
rect -4618 465938 -4534 466174
rect -4298 465938 -4266 466174
rect -4886 465854 -4266 465938
rect -4886 465618 -4854 465854
rect -4618 465618 -4534 465854
rect -4298 465618 -4266 465854
rect -4886 426174 -4266 465618
rect -4886 425938 -4854 426174
rect -4618 425938 -4534 426174
rect -4298 425938 -4266 426174
rect -4886 425854 -4266 425938
rect -4886 425618 -4854 425854
rect -4618 425618 -4534 425854
rect -4298 425618 -4266 425854
rect -4886 386174 -4266 425618
rect -4886 385938 -4854 386174
rect -4618 385938 -4534 386174
rect -4298 385938 -4266 386174
rect -4886 385854 -4266 385938
rect -4886 385618 -4854 385854
rect -4618 385618 -4534 385854
rect -4298 385618 -4266 385854
rect -4886 346174 -4266 385618
rect -4886 345938 -4854 346174
rect -4618 345938 -4534 346174
rect -4298 345938 -4266 346174
rect -4886 345854 -4266 345938
rect -4886 345618 -4854 345854
rect -4618 345618 -4534 345854
rect -4298 345618 -4266 345854
rect -4886 306174 -4266 345618
rect -4886 305938 -4854 306174
rect -4618 305938 -4534 306174
rect -4298 305938 -4266 306174
rect -4886 305854 -4266 305938
rect -4886 305618 -4854 305854
rect -4618 305618 -4534 305854
rect -4298 305618 -4266 305854
rect -4886 266174 -4266 305618
rect -4886 265938 -4854 266174
rect -4618 265938 -4534 266174
rect -4298 265938 -4266 266174
rect -4886 265854 -4266 265938
rect -4886 265618 -4854 265854
rect -4618 265618 -4534 265854
rect -4298 265618 -4266 265854
rect -4886 226174 -4266 265618
rect -4886 225938 -4854 226174
rect -4618 225938 -4534 226174
rect -4298 225938 -4266 226174
rect -4886 225854 -4266 225938
rect -4886 225618 -4854 225854
rect -4618 225618 -4534 225854
rect -4298 225618 -4266 225854
rect -4886 186174 -4266 225618
rect -4886 185938 -4854 186174
rect -4618 185938 -4534 186174
rect -4298 185938 -4266 186174
rect -4886 185854 -4266 185938
rect -4886 185618 -4854 185854
rect -4618 185618 -4534 185854
rect -4298 185618 -4266 185854
rect -4886 146174 -4266 185618
rect -4886 145938 -4854 146174
rect -4618 145938 -4534 146174
rect -4298 145938 -4266 146174
rect -4886 145854 -4266 145938
rect -4886 145618 -4854 145854
rect -4618 145618 -4534 145854
rect -4298 145618 -4266 145854
rect -4886 106174 -4266 145618
rect -4886 105938 -4854 106174
rect -4618 105938 -4534 106174
rect -4298 105938 -4266 106174
rect -4886 105854 -4266 105938
rect -4886 105618 -4854 105854
rect -4618 105618 -4534 105854
rect -4298 105618 -4266 105854
rect -4886 66174 -4266 105618
rect -4886 65938 -4854 66174
rect -4618 65938 -4534 66174
rect -4298 65938 -4266 66174
rect -4886 65854 -4266 65938
rect -4886 65618 -4854 65854
rect -4618 65618 -4534 65854
rect -4298 65618 -4266 65854
rect -4886 26174 -4266 65618
rect -4886 25938 -4854 26174
rect -4618 25938 -4534 26174
rect -4298 25938 -4266 26174
rect -4886 25854 -4266 25938
rect -4886 25618 -4854 25854
rect -4618 25618 -4534 25854
rect -4298 25618 -4266 25854
rect -4886 -3226 -4266 25618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 686174 -3306 706202
rect 4514 706758 5134 707750
rect 4514 706522 4546 706758
rect 4782 706522 4866 706758
rect 5102 706522 5134 706758
rect 4514 706438 5134 706522
rect 4514 706202 4546 706438
rect 4782 706202 4866 706438
rect 5102 706202 5134 706438
rect -3926 685938 -3894 686174
rect -3658 685938 -3574 686174
rect -3338 685938 -3306 686174
rect -3926 685854 -3306 685938
rect -3926 685618 -3894 685854
rect -3658 685618 -3574 685854
rect -3338 685618 -3306 685854
rect -3926 646174 -3306 685618
rect -3926 645938 -3894 646174
rect -3658 645938 -3574 646174
rect -3338 645938 -3306 646174
rect -3926 645854 -3306 645938
rect -3926 645618 -3894 645854
rect -3658 645618 -3574 645854
rect -3338 645618 -3306 645854
rect -3926 606174 -3306 645618
rect -3926 605938 -3894 606174
rect -3658 605938 -3574 606174
rect -3338 605938 -3306 606174
rect -3926 605854 -3306 605938
rect -3926 605618 -3894 605854
rect -3658 605618 -3574 605854
rect -3338 605618 -3306 605854
rect -3926 566174 -3306 605618
rect -3926 565938 -3894 566174
rect -3658 565938 -3574 566174
rect -3338 565938 -3306 566174
rect -3926 565854 -3306 565938
rect -3926 565618 -3894 565854
rect -3658 565618 -3574 565854
rect -3338 565618 -3306 565854
rect -3926 526174 -3306 565618
rect -3926 525938 -3894 526174
rect -3658 525938 -3574 526174
rect -3338 525938 -3306 526174
rect -3926 525854 -3306 525938
rect -3926 525618 -3894 525854
rect -3658 525618 -3574 525854
rect -3338 525618 -3306 525854
rect -3926 486174 -3306 525618
rect -3926 485938 -3894 486174
rect -3658 485938 -3574 486174
rect -3338 485938 -3306 486174
rect -3926 485854 -3306 485938
rect -3926 485618 -3894 485854
rect -3658 485618 -3574 485854
rect -3338 485618 -3306 485854
rect -3926 446174 -3306 485618
rect -3926 445938 -3894 446174
rect -3658 445938 -3574 446174
rect -3338 445938 -3306 446174
rect -3926 445854 -3306 445938
rect -3926 445618 -3894 445854
rect -3658 445618 -3574 445854
rect -3338 445618 -3306 445854
rect -3926 406174 -3306 445618
rect -3926 405938 -3894 406174
rect -3658 405938 -3574 406174
rect -3338 405938 -3306 406174
rect -3926 405854 -3306 405938
rect -3926 405618 -3894 405854
rect -3658 405618 -3574 405854
rect -3338 405618 -3306 405854
rect -3926 366174 -3306 405618
rect -3926 365938 -3894 366174
rect -3658 365938 -3574 366174
rect -3338 365938 -3306 366174
rect -3926 365854 -3306 365938
rect -3926 365618 -3894 365854
rect -3658 365618 -3574 365854
rect -3338 365618 -3306 365854
rect -3926 326174 -3306 365618
rect -3926 325938 -3894 326174
rect -3658 325938 -3574 326174
rect -3338 325938 -3306 326174
rect -3926 325854 -3306 325938
rect -3926 325618 -3894 325854
rect -3658 325618 -3574 325854
rect -3338 325618 -3306 325854
rect -3926 286174 -3306 325618
rect -3926 285938 -3894 286174
rect -3658 285938 -3574 286174
rect -3338 285938 -3306 286174
rect -3926 285854 -3306 285938
rect -3926 285618 -3894 285854
rect -3658 285618 -3574 285854
rect -3338 285618 -3306 285854
rect -3926 246174 -3306 285618
rect -3926 245938 -3894 246174
rect -3658 245938 -3574 246174
rect -3338 245938 -3306 246174
rect -3926 245854 -3306 245938
rect -3926 245618 -3894 245854
rect -3658 245618 -3574 245854
rect -3338 245618 -3306 245854
rect -3926 206174 -3306 245618
rect -3926 205938 -3894 206174
rect -3658 205938 -3574 206174
rect -3338 205938 -3306 206174
rect -3926 205854 -3306 205938
rect -3926 205618 -3894 205854
rect -3658 205618 -3574 205854
rect -3338 205618 -3306 205854
rect -3926 166174 -3306 205618
rect -3926 165938 -3894 166174
rect -3658 165938 -3574 166174
rect -3338 165938 -3306 166174
rect -3926 165854 -3306 165938
rect -3926 165618 -3894 165854
rect -3658 165618 -3574 165854
rect -3338 165618 -3306 165854
rect -3926 126174 -3306 165618
rect -3926 125938 -3894 126174
rect -3658 125938 -3574 126174
rect -3338 125938 -3306 126174
rect -3926 125854 -3306 125938
rect -3926 125618 -3894 125854
rect -3658 125618 -3574 125854
rect -3338 125618 -3306 125854
rect -3926 86174 -3306 125618
rect -3926 85938 -3894 86174
rect -3658 85938 -3574 86174
rect -3338 85938 -3306 86174
rect -3926 85854 -3306 85938
rect -3926 85618 -3894 85854
rect -3658 85618 -3574 85854
rect -3338 85618 -3306 85854
rect -3926 46174 -3306 85618
rect -3926 45938 -3894 46174
rect -3658 45938 -3574 46174
rect -3338 45938 -3306 46174
rect -3926 45854 -3306 45938
rect -3926 45618 -3894 45854
rect -3658 45618 -3574 45854
rect -3338 45618 -3306 45854
rect -3926 6174 -3306 45618
rect -3926 5938 -3894 6174
rect -3658 5938 -3574 6174
rect -3338 5938 -3306 6174
rect -3926 5854 -3306 5938
rect -3926 5618 -3894 5854
rect -3658 5618 -3574 5854
rect -3338 5618 -3306 5854
rect -3926 -2266 -3306 5618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 662454 -2346 705242
rect -2966 662218 -2934 662454
rect -2698 662218 -2614 662454
rect -2378 662218 -2346 662454
rect -2966 662134 -2346 662218
rect -2966 661898 -2934 662134
rect -2698 661898 -2614 662134
rect -2378 661898 -2346 662134
rect -2966 622454 -2346 661898
rect -2966 622218 -2934 622454
rect -2698 622218 -2614 622454
rect -2378 622218 -2346 622454
rect -2966 622134 -2346 622218
rect -2966 621898 -2934 622134
rect -2698 621898 -2614 622134
rect -2378 621898 -2346 622134
rect -2966 582454 -2346 621898
rect -2966 582218 -2934 582454
rect -2698 582218 -2614 582454
rect -2378 582218 -2346 582454
rect -2966 582134 -2346 582218
rect -2966 581898 -2934 582134
rect -2698 581898 -2614 582134
rect -2378 581898 -2346 582134
rect -2966 542454 -2346 581898
rect -2966 542218 -2934 542454
rect -2698 542218 -2614 542454
rect -2378 542218 -2346 542454
rect -2966 542134 -2346 542218
rect -2966 541898 -2934 542134
rect -2698 541898 -2614 542134
rect -2378 541898 -2346 542134
rect -2966 502454 -2346 541898
rect -2966 502218 -2934 502454
rect -2698 502218 -2614 502454
rect -2378 502218 -2346 502454
rect -2966 502134 -2346 502218
rect -2966 501898 -2934 502134
rect -2698 501898 -2614 502134
rect -2378 501898 -2346 502134
rect -2966 462454 -2346 501898
rect -2966 462218 -2934 462454
rect -2698 462218 -2614 462454
rect -2378 462218 -2346 462454
rect -2966 462134 -2346 462218
rect -2966 461898 -2934 462134
rect -2698 461898 -2614 462134
rect -2378 461898 -2346 462134
rect -2966 422454 -2346 461898
rect -2966 422218 -2934 422454
rect -2698 422218 -2614 422454
rect -2378 422218 -2346 422454
rect -2966 422134 -2346 422218
rect -2966 421898 -2934 422134
rect -2698 421898 -2614 422134
rect -2378 421898 -2346 422134
rect -2966 382454 -2346 421898
rect -2966 382218 -2934 382454
rect -2698 382218 -2614 382454
rect -2378 382218 -2346 382454
rect -2966 382134 -2346 382218
rect -2966 381898 -2934 382134
rect -2698 381898 -2614 382134
rect -2378 381898 -2346 382134
rect -2966 342454 -2346 381898
rect -2966 342218 -2934 342454
rect -2698 342218 -2614 342454
rect -2378 342218 -2346 342454
rect -2966 342134 -2346 342218
rect -2966 341898 -2934 342134
rect -2698 341898 -2614 342134
rect -2378 341898 -2346 342134
rect -2966 302454 -2346 341898
rect -2966 302218 -2934 302454
rect -2698 302218 -2614 302454
rect -2378 302218 -2346 302454
rect -2966 302134 -2346 302218
rect -2966 301898 -2934 302134
rect -2698 301898 -2614 302134
rect -2378 301898 -2346 302134
rect -2966 262454 -2346 301898
rect -2966 262218 -2934 262454
rect -2698 262218 -2614 262454
rect -2378 262218 -2346 262454
rect -2966 262134 -2346 262218
rect -2966 261898 -2934 262134
rect -2698 261898 -2614 262134
rect -2378 261898 -2346 262134
rect -2966 222454 -2346 261898
rect -2966 222218 -2934 222454
rect -2698 222218 -2614 222454
rect -2378 222218 -2346 222454
rect -2966 222134 -2346 222218
rect -2966 221898 -2934 222134
rect -2698 221898 -2614 222134
rect -2378 221898 -2346 222134
rect -2966 182454 -2346 221898
rect -2966 182218 -2934 182454
rect -2698 182218 -2614 182454
rect -2378 182218 -2346 182454
rect -2966 182134 -2346 182218
rect -2966 181898 -2934 182134
rect -2698 181898 -2614 182134
rect -2378 181898 -2346 182134
rect -2966 142454 -2346 181898
rect -2966 142218 -2934 142454
rect -2698 142218 -2614 142454
rect -2378 142218 -2346 142454
rect -2966 142134 -2346 142218
rect -2966 141898 -2934 142134
rect -2698 141898 -2614 142134
rect -2378 141898 -2346 142134
rect -2966 102454 -2346 141898
rect -2966 102218 -2934 102454
rect -2698 102218 -2614 102454
rect -2378 102218 -2346 102454
rect -2966 102134 -2346 102218
rect -2966 101898 -2934 102134
rect -2698 101898 -2614 102134
rect -2378 101898 -2346 102134
rect -2966 62454 -2346 101898
rect -2966 62218 -2934 62454
rect -2698 62218 -2614 62454
rect -2378 62218 -2346 62454
rect -2966 62134 -2346 62218
rect -2966 61898 -2934 62134
rect -2698 61898 -2614 62134
rect -2378 61898 -2346 62134
rect -2966 22454 -2346 61898
rect -2966 22218 -2934 22454
rect -2698 22218 -2614 22454
rect -2378 22218 -2346 22454
rect -2966 22134 -2346 22218
rect -2966 21898 -2934 22134
rect -2698 21898 -2614 22134
rect -2378 21898 -2346 22134
rect -2966 -1306 -2346 21898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 682454 -1386 704282
rect -2006 682218 -1974 682454
rect -1738 682218 -1654 682454
rect -1418 682218 -1386 682454
rect -2006 682134 -1386 682218
rect -2006 681898 -1974 682134
rect -1738 681898 -1654 682134
rect -1418 681898 -1386 682134
rect -2006 642454 -1386 681898
rect -2006 642218 -1974 642454
rect -1738 642218 -1654 642454
rect -1418 642218 -1386 642454
rect -2006 642134 -1386 642218
rect -2006 641898 -1974 642134
rect -1738 641898 -1654 642134
rect -1418 641898 -1386 642134
rect -2006 602454 -1386 641898
rect -2006 602218 -1974 602454
rect -1738 602218 -1654 602454
rect -1418 602218 -1386 602454
rect -2006 602134 -1386 602218
rect -2006 601898 -1974 602134
rect -1738 601898 -1654 602134
rect -1418 601898 -1386 602134
rect -2006 562454 -1386 601898
rect -2006 562218 -1974 562454
rect -1738 562218 -1654 562454
rect -1418 562218 -1386 562454
rect -2006 562134 -1386 562218
rect -2006 561898 -1974 562134
rect -1738 561898 -1654 562134
rect -1418 561898 -1386 562134
rect -2006 522454 -1386 561898
rect -2006 522218 -1974 522454
rect -1738 522218 -1654 522454
rect -1418 522218 -1386 522454
rect -2006 522134 -1386 522218
rect -2006 521898 -1974 522134
rect -1738 521898 -1654 522134
rect -1418 521898 -1386 522134
rect -2006 482454 -1386 521898
rect -2006 482218 -1974 482454
rect -1738 482218 -1654 482454
rect -1418 482218 -1386 482454
rect -2006 482134 -1386 482218
rect -2006 481898 -1974 482134
rect -1738 481898 -1654 482134
rect -1418 481898 -1386 482134
rect -2006 442454 -1386 481898
rect -2006 442218 -1974 442454
rect -1738 442218 -1654 442454
rect -1418 442218 -1386 442454
rect -2006 442134 -1386 442218
rect -2006 441898 -1974 442134
rect -1738 441898 -1654 442134
rect -1418 441898 -1386 442134
rect -2006 402454 -1386 441898
rect -2006 402218 -1974 402454
rect -1738 402218 -1654 402454
rect -1418 402218 -1386 402454
rect -2006 402134 -1386 402218
rect -2006 401898 -1974 402134
rect -1738 401898 -1654 402134
rect -1418 401898 -1386 402134
rect -2006 362454 -1386 401898
rect -2006 362218 -1974 362454
rect -1738 362218 -1654 362454
rect -1418 362218 -1386 362454
rect -2006 362134 -1386 362218
rect -2006 361898 -1974 362134
rect -1738 361898 -1654 362134
rect -1418 361898 -1386 362134
rect -2006 322454 -1386 361898
rect -2006 322218 -1974 322454
rect -1738 322218 -1654 322454
rect -1418 322218 -1386 322454
rect -2006 322134 -1386 322218
rect -2006 321898 -1974 322134
rect -1738 321898 -1654 322134
rect -1418 321898 -1386 322134
rect -2006 282454 -1386 321898
rect -2006 282218 -1974 282454
rect -1738 282218 -1654 282454
rect -1418 282218 -1386 282454
rect -2006 282134 -1386 282218
rect -2006 281898 -1974 282134
rect -1738 281898 -1654 282134
rect -1418 281898 -1386 282134
rect -2006 242454 -1386 281898
rect -2006 242218 -1974 242454
rect -1738 242218 -1654 242454
rect -1418 242218 -1386 242454
rect -2006 242134 -1386 242218
rect -2006 241898 -1974 242134
rect -1738 241898 -1654 242134
rect -1418 241898 -1386 242134
rect -2006 202454 -1386 241898
rect -2006 202218 -1974 202454
rect -1738 202218 -1654 202454
rect -1418 202218 -1386 202454
rect -2006 202134 -1386 202218
rect -2006 201898 -1974 202134
rect -1738 201898 -1654 202134
rect -1418 201898 -1386 202134
rect -2006 162454 -1386 201898
rect -2006 162218 -1974 162454
rect -1738 162218 -1654 162454
rect -1418 162218 -1386 162454
rect -2006 162134 -1386 162218
rect -2006 161898 -1974 162134
rect -1738 161898 -1654 162134
rect -1418 161898 -1386 162134
rect -2006 122454 -1386 161898
rect -2006 122218 -1974 122454
rect -1738 122218 -1654 122454
rect -1418 122218 -1386 122454
rect -2006 122134 -1386 122218
rect -2006 121898 -1974 122134
rect -1738 121898 -1654 122134
rect -1418 121898 -1386 122134
rect -2006 82454 -1386 121898
rect -2006 82218 -1974 82454
rect -1738 82218 -1654 82454
rect -1418 82218 -1386 82454
rect -2006 82134 -1386 82218
rect -2006 81898 -1974 82134
rect -1738 81898 -1654 82134
rect -1418 81898 -1386 82134
rect -2006 42454 -1386 81898
rect -2006 42218 -1974 42454
rect -1738 42218 -1654 42454
rect -1418 42218 -1386 42454
rect -2006 42134 -1386 42218
rect -2006 41898 -1974 42134
rect -1738 41898 -1654 42134
rect -1418 41898 -1386 42134
rect -2006 2454 -1386 41898
rect -2006 2218 -1974 2454
rect -1738 2218 -1654 2454
rect -1418 2218 -1386 2454
rect -2006 2134 -1386 2218
rect -2006 1898 -1974 2134
rect -1738 1898 -1654 2134
rect -1418 1898 -1386 2134
rect -2006 -346 -1386 1898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 794 704838 1414 705830
rect 794 704602 826 704838
rect 1062 704602 1146 704838
rect 1382 704602 1414 704838
rect 794 704518 1414 704602
rect 794 704282 826 704518
rect 1062 704282 1146 704518
rect 1382 704282 1414 704518
rect 794 682454 1414 704282
rect 794 682218 826 682454
rect 1062 682218 1146 682454
rect 1382 682218 1414 682454
rect 794 682134 1414 682218
rect 794 681898 826 682134
rect 1062 681898 1146 682134
rect 1382 681898 1414 682134
rect 794 642454 1414 681898
rect 794 642218 826 642454
rect 1062 642218 1146 642454
rect 1382 642218 1414 642454
rect 794 642134 1414 642218
rect 794 641898 826 642134
rect 1062 641898 1146 642134
rect 1382 641898 1414 642134
rect 794 602454 1414 641898
rect 794 602218 826 602454
rect 1062 602218 1146 602454
rect 1382 602218 1414 602454
rect 794 602134 1414 602218
rect 794 601898 826 602134
rect 1062 601898 1146 602134
rect 1382 601898 1414 602134
rect 794 562454 1414 601898
rect 794 562218 826 562454
rect 1062 562218 1146 562454
rect 1382 562218 1414 562454
rect 794 562134 1414 562218
rect 794 561898 826 562134
rect 1062 561898 1146 562134
rect 1382 561898 1414 562134
rect 794 522454 1414 561898
rect 794 522218 826 522454
rect 1062 522218 1146 522454
rect 1382 522218 1414 522454
rect 794 522134 1414 522218
rect 794 521898 826 522134
rect 1062 521898 1146 522134
rect 1382 521898 1414 522134
rect 794 482454 1414 521898
rect 794 482218 826 482454
rect 1062 482218 1146 482454
rect 1382 482218 1414 482454
rect 794 482134 1414 482218
rect 794 481898 826 482134
rect 1062 481898 1146 482134
rect 1382 481898 1414 482134
rect 794 442454 1414 481898
rect 794 442218 826 442454
rect 1062 442218 1146 442454
rect 1382 442218 1414 442454
rect 794 442134 1414 442218
rect 794 441898 826 442134
rect 1062 441898 1146 442134
rect 1382 441898 1414 442134
rect 794 402454 1414 441898
rect 794 402218 826 402454
rect 1062 402218 1146 402454
rect 1382 402218 1414 402454
rect 794 402134 1414 402218
rect 794 401898 826 402134
rect 1062 401898 1146 402134
rect 1382 401898 1414 402134
rect 794 362454 1414 401898
rect 794 362218 826 362454
rect 1062 362218 1146 362454
rect 1382 362218 1414 362454
rect 794 362134 1414 362218
rect 794 361898 826 362134
rect 1062 361898 1146 362134
rect 1382 361898 1414 362134
rect 794 322454 1414 361898
rect 794 322218 826 322454
rect 1062 322218 1146 322454
rect 1382 322218 1414 322454
rect 794 322134 1414 322218
rect 794 321898 826 322134
rect 1062 321898 1146 322134
rect 1382 321898 1414 322134
rect 794 282454 1414 321898
rect 794 282218 826 282454
rect 1062 282218 1146 282454
rect 1382 282218 1414 282454
rect 794 282134 1414 282218
rect 794 281898 826 282134
rect 1062 281898 1146 282134
rect 1382 281898 1414 282134
rect 794 242454 1414 281898
rect 794 242218 826 242454
rect 1062 242218 1146 242454
rect 1382 242218 1414 242454
rect 794 242134 1414 242218
rect 794 241898 826 242134
rect 1062 241898 1146 242134
rect 1382 241898 1414 242134
rect 794 202454 1414 241898
rect 794 202218 826 202454
rect 1062 202218 1146 202454
rect 1382 202218 1414 202454
rect 794 202134 1414 202218
rect 794 201898 826 202134
rect 1062 201898 1146 202134
rect 1382 201898 1414 202134
rect 794 162454 1414 201898
rect 794 162218 826 162454
rect 1062 162218 1146 162454
rect 1382 162218 1414 162454
rect 794 162134 1414 162218
rect 794 161898 826 162134
rect 1062 161898 1146 162134
rect 1382 161898 1414 162134
rect 794 122454 1414 161898
rect 794 122218 826 122454
rect 1062 122218 1146 122454
rect 1382 122218 1414 122454
rect 794 122134 1414 122218
rect 794 121898 826 122134
rect 1062 121898 1146 122134
rect 1382 121898 1414 122134
rect 794 82454 1414 121898
rect 794 82218 826 82454
rect 1062 82218 1146 82454
rect 1382 82218 1414 82454
rect 794 82134 1414 82218
rect 794 81898 826 82134
rect 1062 81898 1146 82134
rect 1382 81898 1414 82134
rect 794 42454 1414 81898
rect 794 42218 826 42454
rect 1062 42218 1146 42454
rect 1382 42218 1414 42454
rect 794 42134 1414 42218
rect 794 41898 826 42134
rect 1062 41898 1146 42134
rect 1382 41898 1414 42134
rect 794 2454 1414 41898
rect 794 2218 826 2454
rect 1062 2218 1146 2454
rect 1382 2218 1414 2454
rect 794 2134 1414 2218
rect 794 1898 826 2134
rect 1062 1898 1146 2134
rect 1382 1898 1414 2134
rect 794 -346 1414 1898
rect 794 -582 826 -346
rect 1062 -582 1146 -346
rect 1382 -582 1414 -346
rect 794 -666 1414 -582
rect 794 -902 826 -666
rect 1062 -902 1146 -666
rect 1382 -902 1414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 794 -1894 1414 -902
rect 4514 686174 5134 706202
rect 4514 685938 4546 686174
rect 4782 685938 4866 686174
rect 5102 685938 5134 686174
rect 4514 685854 5134 685938
rect 4514 685618 4546 685854
rect 4782 685618 4866 685854
rect 5102 685618 5134 685854
rect 4514 646174 5134 685618
rect 4514 645938 4546 646174
rect 4782 645938 4866 646174
rect 5102 645938 5134 646174
rect 4514 645854 5134 645938
rect 4514 645618 4546 645854
rect 4782 645618 4866 645854
rect 5102 645618 5134 645854
rect 4514 606174 5134 645618
rect 4514 605938 4546 606174
rect 4782 605938 4866 606174
rect 5102 605938 5134 606174
rect 4514 605854 5134 605938
rect 4514 605618 4546 605854
rect 4782 605618 4866 605854
rect 5102 605618 5134 605854
rect 4514 566174 5134 605618
rect 4514 565938 4546 566174
rect 4782 565938 4866 566174
rect 5102 565938 5134 566174
rect 4514 565854 5134 565938
rect 4514 565618 4546 565854
rect 4782 565618 4866 565854
rect 5102 565618 5134 565854
rect 4514 526174 5134 565618
rect 4514 525938 4546 526174
rect 4782 525938 4866 526174
rect 5102 525938 5134 526174
rect 4514 525854 5134 525938
rect 4514 525618 4546 525854
rect 4782 525618 4866 525854
rect 5102 525618 5134 525854
rect 4514 486174 5134 525618
rect 4514 485938 4546 486174
rect 4782 485938 4866 486174
rect 5102 485938 5134 486174
rect 4514 485854 5134 485938
rect 4514 485618 4546 485854
rect 4782 485618 4866 485854
rect 5102 485618 5134 485854
rect 4514 446174 5134 485618
rect 4514 445938 4546 446174
rect 4782 445938 4866 446174
rect 5102 445938 5134 446174
rect 4514 445854 5134 445938
rect 4514 445618 4546 445854
rect 4782 445618 4866 445854
rect 5102 445618 5134 445854
rect 4514 406174 5134 445618
rect 4514 405938 4546 406174
rect 4782 405938 4866 406174
rect 5102 405938 5134 406174
rect 4514 405854 5134 405938
rect 4514 405618 4546 405854
rect 4782 405618 4866 405854
rect 5102 405618 5134 405854
rect 4514 366174 5134 405618
rect 4514 365938 4546 366174
rect 4782 365938 4866 366174
rect 5102 365938 5134 366174
rect 4514 365854 5134 365938
rect 4514 365618 4546 365854
rect 4782 365618 4866 365854
rect 5102 365618 5134 365854
rect 4514 326174 5134 365618
rect 4514 325938 4546 326174
rect 4782 325938 4866 326174
rect 5102 325938 5134 326174
rect 4514 325854 5134 325938
rect 4514 325618 4546 325854
rect 4782 325618 4866 325854
rect 5102 325618 5134 325854
rect 4514 286174 5134 325618
rect 4514 285938 4546 286174
rect 4782 285938 4866 286174
rect 5102 285938 5134 286174
rect 4514 285854 5134 285938
rect 4514 285618 4546 285854
rect 4782 285618 4866 285854
rect 5102 285618 5134 285854
rect 4514 246174 5134 285618
rect 4514 245938 4546 246174
rect 4782 245938 4866 246174
rect 5102 245938 5134 246174
rect 4514 245854 5134 245938
rect 4514 245618 4546 245854
rect 4782 245618 4866 245854
rect 5102 245618 5134 245854
rect 4514 206174 5134 245618
rect 4514 205938 4546 206174
rect 4782 205938 4866 206174
rect 5102 205938 5134 206174
rect 4514 205854 5134 205938
rect 4514 205618 4546 205854
rect 4782 205618 4866 205854
rect 5102 205618 5134 205854
rect 4514 166174 5134 205618
rect 4514 165938 4546 166174
rect 4782 165938 4866 166174
rect 5102 165938 5134 166174
rect 4514 165854 5134 165938
rect 4514 165618 4546 165854
rect 4782 165618 4866 165854
rect 5102 165618 5134 165854
rect 4514 126174 5134 165618
rect 4514 125938 4546 126174
rect 4782 125938 4866 126174
rect 5102 125938 5134 126174
rect 4514 125854 5134 125938
rect 4514 125618 4546 125854
rect 4782 125618 4866 125854
rect 5102 125618 5134 125854
rect 4514 86174 5134 125618
rect 4514 85938 4546 86174
rect 4782 85938 4866 86174
rect 5102 85938 5134 86174
rect 4514 85854 5134 85938
rect 4514 85618 4546 85854
rect 4782 85618 4866 85854
rect 5102 85618 5134 85854
rect 4514 46174 5134 85618
rect 4514 45938 4546 46174
rect 4782 45938 4866 46174
rect 5102 45938 5134 46174
rect 4514 45854 5134 45938
rect 4514 45618 4546 45854
rect 4782 45618 4866 45854
rect 5102 45618 5134 45854
rect 4514 6174 5134 45618
rect 4514 5938 4546 6174
rect 4782 5938 4866 6174
rect 5102 5938 5134 6174
rect 4514 5854 5134 5938
rect 4514 5618 4546 5854
rect 4782 5618 4866 5854
rect 5102 5618 5134 5854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 4514 -2266 5134 5618
rect 4514 -2502 4546 -2266
rect 4782 -2502 4866 -2266
rect 5102 -2502 5134 -2266
rect 4514 -2586 5134 -2502
rect 4514 -2822 4546 -2586
rect 4782 -2822 4866 -2586
rect 5102 -2822 5134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 4514 -3814 5134 -2822
rect 8234 689894 8854 708122
rect 8234 689658 8266 689894
rect 8502 689658 8586 689894
rect 8822 689658 8854 689894
rect 8234 689574 8854 689658
rect 8234 689338 8266 689574
rect 8502 689338 8586 689574
rect 8822 689338 8854 689574
rect 8234 649894 8854 689338
rect 8234 649658 8266 649894
rect 8502 649658 8586 649894
rect 8822 649658 8854 649894
rect 8234 649574 8854 649658
rect 8234 649338 8266 649574
rect 8502 649338 8586 649574
rect 8822 649338 8854 649574
rect 8234 609894 8854 649338
rect 8234 609658 8266 609894
rect 8502 609658 8586 609894
rect 8822 609658 8854 609894
rect 8234 609574 8854 609658
rect 8234 609338 8266 609574
rect 8502 609338 8586 609574
rect 8822 609338 8854 609574
rect 8234 569894 8854 609338
rect 8234 569658 8266 569894
rect 8502 569658 8586 569894
rect 8822 569658 8854 569894
rect 8234 569574 8854 569658
rect 8234 569338 8266 569574
rect 8502 569338 8586 569574
rect 8822 569338 8854 569574
rect 8234 529894 8854 569338
rect 8234 529658 8266 529894
rect 8502 529658 8586 529894
rect 8822 529658 8854 529894
rect 8234 529574 8854 529658
rect 8234 529338 8266 529574
rect 8502 529338 8586 529574
rect 8822 529338 8854 529574
rect 8234 489894 8854 529338
rect 8234 489658 8266 489894
rect 8502 489658 8586 489894
rect 8822 489658 8854 489894
rect 8234 489574 8854 489658
rect 8234 489338 8266 489574
rect 8502 489338 8586 489574
rect 8822 489338 8854 489574
rect 8234 449894 8854 489338
rect 8234 449658 8266 449894
rect 8502 449658 8586 449894
rect 8822 449658 8854 449894
rect 8234 449574 8854 449658
rect 8234 449338 8266 449574
rect 8502 449338 8586 449574
rect 8822 449338 8854 449574
rect 8234 409894 8854 449338
rect 8234 409658 8266 409894
rect 8502 409658 8586 409894
rect 8822 409658 8854 409894
rect 8234 409574 8854 409658
rect 8234 409338 8266 409574
rect 8502 409338 8586 409574
rect 8822 409338 8854 409574
rect 8234 369894 8854 409338
rect 8234 369658 8266 369894
rect 8502 369658 8586 369894
rect 8822 369658 8854 369894
rect 8234 369574 8854 369658
rect 8234 369338 8266 369574
rect 8502 369338 8586 369574
rect 8822 369338 8854 369574
rect 8234 329894 8854 369338
rect 8234 329658 8266 329894
rect 8502 329658 8586 329894
rect 8822 329658 8854 329894
rect 8234 329574 8854 329658
rect 8234 329338 8266 329574
rect 8502 329338 8586 329574
rect 8822 329338 8854 329574
rect 8234 289894 8854 329338
rect 8234 289658 8266 289894
rect 8502 289658 8586 289894
rect 8822 289658 8854 289894
rect 8234 289574 8854 289658
rect 8234 289338 8266 289574
rect 8502 289338 8586 289574
rect 8822 289338 8854 289574
rect 8234 249894 8854 289338
rect 8234 249658 8266 249894
rect 8502 249658 8586 249894
rect 8822 249658 8854 249894
rect 8234 249574 8854 249658
rect 8234 249338 8266 249574
rect 8502 249338 8586 249574
rect 8822 249338 8854 249574
rect 8234 209894 8854 249338
rect 8234 209658 8266 209894
rect 8502 209658 8586 209894
rect 8822 209658 8854 209894
rect 8234 209574 8854 209658
rect 8234 209338 8266 209574
rect 8502 209338 8586 209574
rect 8822 209338 8854 209574
rect 8234 169894 8854 209338
rect 8234 169658 8266 169894
rect 8502 169658 8586 169894
rect 8822 169658 8854 169894
rect 8234 169574 8854 169658
rect 8234 169338 8266 169574
rect 8502 169338 8586 169574
rect 8822 169338 8854 169574
rect 8234 129894 8854 169338
rect 8234 129658 8266 129894
rect 8502 129658 8586 129894
rect 8822 129658 8854 129894
rect 8234 129574 8854 129658
rect 8234 129338 8266 129574
rect 8502 129338 8586 129574
rect 8822 129338 8854 129574
rect 8234 89894 8854 129338
rect 8234 89658 8266 89894
rect 8502 89658 8586 89894
rect 8822 89658 8854 89894
rect 8234 89574 8854 89658
rect 8234 89338 8266 89574
rect 8502 89338 8586 89574
rect 8822 89338 8854 89574
rect 8234 49894 8854 89338
rect 8234 49658 8266 49894
rect 8502 49658 8586 49894
rect 8822 49658 8854 49894
rect 8234 49574 8854 49658
rect 8234 49338 8266 49574
rect 8502 49338 8586 49574
rect 8822 49338 8854 49574
rect 8234 9894 8854 49338
rect 8234 9658 8266 9894
rect 8502 9658 8586 9894
rect 8822 9658 8854 9894
rect 8234 9574 8854 9658
rect 8234 9338 8266 9574
rect 8502 9338 8586 9574
rect 8822 9338 8854 9574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 8234 -4186 8854 9338
rect 8234 -4422 8266 -4186
rect 8502 -4422 8586 -4186
rect 8822 -4422 8854 -4186
rect 8234 -4506 8854 -4422
rect 8234 -4742 8266 -4506
rect 8502 -4742 8586 -4506
rect 8822 -4742 8854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 8234 -5734 8854 -4742
rect 11954 693614 12574 710042
rect 31954 711558 32574 711590
rect 31954 711322 31986 711558
rect 32222 711322 32306 711558
rect 32542 711322 32574 711558
rect 31954 711238 32574 711322
rect 31954 711002 31986 711238
rect 32222 711002 32306 711238
rect 32542 711002 32574 711238
rect 28234 709638 28854 709670
rect 28234 709402 28266 709638
rect 28502 709402 28586 709638
rect 28822 709402 28854 709638
rect 28234 709318 28854 709402
rect 28234 709082 28266 709318
rect 28502 709082 28586 709318
rect 28822 709082 28854 709318
rect 24514 707718 25134 707750
rect 24514 707482 24546 707718
rect 24782 707482 24866 707718
rect 25102 707482 25134 707718
rect 24514 707398 25134 707482
rect 24514 707162 24546 707398
rect 24782 707162 24866 707398
rect 25102 707162 25134 707398
rect 11954 693378 11986 693614
rect 12222 693378 12306 693614
rect 12542 693378 12574 693614
rect 11954 693294 12574 693378
rect 11954 693058 11986 693294
rect 12222 693058 12306 693294
rect 12542 693058 12574 693294
rect 11954 653614 12574 693058
rect 11954 653378 11986 653614
rect 12222 653378 12306 653614
rect 12542 653378 12574 653614
rect 11954 653294 12574 653378
rect 11954 653058 11986 653294
rect 12222 653058 12306 653294
rect 12542 653058 12574 653294
rect 11954 613614 12574 653058
rect 11954 613378 11986 613614
rect 12222 613378 12306 613614
rect 12542 613378 12574 613614
rect 11954 613294 12574 613378
rect 11954 613058 11986 613294
rect 12222 613058 12306 613294
rect 12542 613058 12574 613294
rect 11954 573614 12574 613058
rect 11954 573378 11986 573614
rect 12222 573378 12306 573614
rect 12542 573378 12574 573614
rect 11954 573294 12574 573378
rect 11954 573058 11986 573294
rect 12222 573058 12306 573294
rect 12542 573058 12574 573294
rect 11954 533614 12574 573058
rect 11954 533378 11986 533614
rect 12222 533378 12306 533614
rect 12542 533378 12574 533614
rect 11954 533294 12574 533378
rect 11954 533058 11986 533294
rect 12222 533058 12306 533294
rect 12542 533058 12574 533294
rect 11954 493614 12574 533058
rect 11954 493378 11986 493614
rect 12222 493378 12306 493614
rect 12542 493378 12574 493614
rect 11954 493294 12574 493378
rect 11954 493058 11986 493294
rect 12222 493058 12306 493294
rect 12542 493058 12574 493294
rect 11954 453614 12574 493058
rect 11954 453378 11986 453614
rect 12222 453378 12306 453614
rect 12542 453378 12574 453614
rect 11954 453294 12574 453378
rect 11954 453058 11986 453294
rect 12222 453058 12306 453294
rect 12542 453058 12574 453294
rect 11954 413614 12574 453058
rect 11954 413378 11986 413614
rect 12222 413378 12306 413614
rect 12542 413378 12574 413614
rect 11954 413294 12574 413378
rect 11954 413058 11986 413294
rect 12222 413058 12306 413294
rect 12542 413058 12574 413294
rect 11954 373614 12574 413058
rect 11954 373378 11986 373614
rect 12222 373378 12306 373614
rect 12542 373378 12574 373614
rect 11954 373294 12574 373378
rect 11954 373058 11986 373294
rect 12222 373058 12306 373294
rect 12542 373058 12574 373294
rect 11954 333614 12574 373058
rect 11954 333378 11986 333614
rect 12222 333378 12306 333614
rect 12542 333378 12574 333614
rect 11954 333294 12574 333378
rect 11954 333058 11986 333294
rect 12222 333058 12306 333294
rect 12542 333058 12574 333294
rect 11954 293614 12574 333058
rect 11954 293378 11986 293614
rect 12222 293378 12306 293614
rect 12542 293378 12574 293614
rect 11954 293294 12574 293378
rect 11954 293058 11986 293294
rect 12222 293058 12306 293294
rect 12542 293058 12574 293294
rect 11954 253614 12574 293058
rect 11954 253378 11986 253614
rect 12222 253378 12306 253614
rect 12542 253378 12574 253614
rect 11954 253294 12574 253378
rect 11954 253058 11986 253294
rect 12222 253058 12306 253294
rect 12542 253058 12574 253294
rect 11954 213614 12574 253058
rect 11954 213378 11986 213614
rect 12222 213378 12306 213614
rect 12542 213378 12574 213614
rect 11954 213294 12574 213378
rect 11954 213058 11986 213294
rect 12222 213058 12306 213294
rect 12542 213058 12574 213294
rect 11954 173614 12574 213058
rect 11954 173378 11986 173614
rect 12222 173378 12306 173614
rect 12542 173378 12574 173614
rect 11954 173294 12574 173378
rect 11954 173058 11986 173294
rect 12222 173058 12306 173294
rect 12542 173058 12574 173294
rect 11954 133614 12574 173058
rect 11954 133378 11986 133614
rect 12222 133378 12306 133614
rect 12542 133378 12574 133614
rect 11954 133294 12574 133378
rect 11954 133058 11986 133294
rect 12222 133058 12306 133294
rect 12542 133058 12574 133294
rect 11954 93614 12574 133058
rect 11954 93378 11986 93614
rect 12222 93378 12306 93614
rect 12542 93378 12574 93614
rect 11954 93294 12574 93378
rect 11954 93058 11986 93294
rect 12222 93058 12306 93294
rect 12542 93058 12574 93294
rect 11954 53614 12574 93058
rect 11954 53378 11986 53614
rect 12222 53378 12306 53614
rect 12542 53378 12574 53614
rect 11954 53294 12574 53378
rect 11954 53058 11986 53294
rect 12222 53058 12306 53294
rect 12542 53058 12574 53294
rect 11954 13614 12574 53058
rect 11954 13378 11986 13614
rect 12222 13378 12306 13614
rect 12542 13378 12574 13614
rect 11954 13294 12574 13378
rect 11954 13058 11986 13294
rect 12222 13058 12306 13294
rect 12542 13058 12574 13294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 11954 -6106 12574 13058
rect 20794 705798 21414 705830
rect 20794 705562 20826 705798
rect 21062 705562 21146 705798
rect 21382 705562 21414 705798
rect 20794 705478 21414 705562
rect 20794 705242 20826 705478
rect 21062 705242 21146 705478
rect 21382 705242 21414 705478
rect 20794 662454 21414 705242
rect 20794 662218 20826 662454
rect 21062 662218 21146 662454
rect 21382 662218 21414 662454
rect 20794 662134 21414 662218
rect 20794 661898 20826 662134
rect 21062 661898 21146 662134
rect 21382 661898 21414 662134
rect 20794 622454 21414 661898
rect 20794 622218 20826 622454
rect 21062 622218 21146 622454
rect 21382 622218 21414 622454
rect 20794 622134 21414 622218
rect 20794 621898 20826 622134
rect 21062 621898 21146 622134
rect 21382 621898 21414 622134
rect 20794 582454 21414 621898
rect 20794 582218 20826 582454
rect 21062 582218 21146 582454
rect 21382 582218 21414 582454
rect 20794 582134 21414 582218
rect 20794 581898 20826 582134
rect 21062 581898 21146 582134
rect 21382 581898 21414 582134
rect 20794 542454 21414 581898
rect 20794 542218 20826 542454
rect 21062 542218 21146 542454
rect 21382 542218 21414 542454
rect 20794 542134 21414 542218
rect 20794 541898 20826 542134
rect 21062 541898 21146 542134
rect 21382 541898 21414 542134
rect 20794 502454 21414 541898
rect 20794 502218 20826 502454
rect 21062 502218 21146 502454
rect 21382 502218 21414 502454
rect 20794 502134 21414 502218
rect 20794 501898 20826 502134
rect 21062 501898 21146 502134
rect 21382 501898 21414 502134
rect 20794 462454 21414 501898
rect 20794 462218 20826 462454
rect 21062 462218 21146 462454
rect 21382 462218 21414 462454
rect 20794 462134 21414 462218
rect 20794 461898 20826 462134
rect 21062 461898 21146 462134
rect 21382 461898 21414 462134
rect 20794 422454 21414 461898
rect 20794 422218 20826 422454
rect 21062 422218 21146 422454
rect 21382 422218 21414 422454
rect 20794 422134 21414 422218
rect 20794 421898 20826 422134
rect 21062 421898 21146 422134
rect 21382 421898 21414 422134
rect 20794 382454 21414 421898
rect 20794 382218 20826 382454
rect 21062 382218 21146 382454
rect 21382 382218 21414 382454
rect 20794 382134 21414 382218
rect 20794 381898 20826 382134
rect 21062 381898 21146 382134
rect 21382 381898 21414 382134
rect 20794 342454 21414 381898
rect 20794 342218 20826 342454
rect 21062 342218 21146 342454
rect 21382 342218 21414 342454
rect 20794 342134 21414 342218
rect 20794 341898 20826 342134
rect 21062 341898 21146 342134
rect 21382 341898 21414 342134
rect 20794 302454 21414 341898
rect 20794 302218 20826 302454
rect 21062 302218 21146 302454
rect 21382 302218 21414 302454
rect 20794 302134 21414 302218
rect 20794 301898 20826 302134
rect 21062 301898 21146 302134
rect 21382 301898 21414 302134
rect 20794 262454 21414 301898
rect 20794 262218 20826 262454
rect 21062 262218 21146 262454
rect 21382 262218 21414 262454
rect 20794 262134 21414 262218
rect 20794 261898 20826 262134
rect 21062 261898 21146 262134
rect 21382 261898 21414 262134
rect 20794 222454 21414 261898
rect 20794 222218 20826 222454
rect 21062 222218 21146 222454
rect 21382 222218 21414 222454
rect 20794 222134 21414 222218
rect 20794 221898 20826 222134
rect 21062 221898 21146 222134
rect 21382 221898 21414 222134
rect 20794 182454 21414 221898
rect 20794 182218 20826 182454
rect 21062 182218 21146 182454
rect 21382 182218 21414 182454
rect 20794 182134 21414 182218
rect 20794 181898 20826 182134
rect 21062 181898 21146 182134
rect 21382 181898 21414 182134
rect 20794 142454 21414 181898
rect 20794 142218 20826 142454
rect 21062 142218 21146 142454
rect 21382 142218 21414 142454
rect 20794 142134 21414 142218
rect 20794 141898 20826 142134
rect 21062 141898 21146 142134
rect 21382 141898 21414 142134
rect 20794 102454 21414 141898
rect 20794 102218 20826 102454
rect 21062 102218 21146 102454
rect 21382 102218 21414 102454
rect 20794 102134 21414 102218
rect 20794 101898 20826 102134
rect 21062 101898 21146 102134
rect 21382 101898 21414 102134
rect 20794 62454 21414 101898
rect 20794 62218 20826 62454
rect 21062 62218 21146 62454
rect 21382 62218 21414 62454
rect 20794 62134 21414 62218
rect 20794 61898 20826 62134
rect 21062 61898 21146 62134
rect 21382 61898 21414 62134
rect 20794 22454 21414 61898
rect 20794 22218 20826 22454
rect 21062 22218 21146 22454
rect 21382 22218 21414 22454
rect 20794 22134 21414 22218
rect 20794 21898 20826 22134
rect 21062 21898 21146 22134
rect 21382 21898 21414 22134
rect 20794 -1306 21414 21898
rect 20794 -1542 20826 -1306
rect 21062 -1542 21146 -1306
rect 21382 -1542 21414 -1306
rect 20794 -1626 21414 -1542
rect 20794 -1862 20826 -1626
rect 21062 -1862 21146 -1626
rect 21382 -1862 21414 -1626
rect 20794 -1894 21414 -1862
rect 24514 666174 25134 707162
rect 24514 665938 24546 666174
rect 24782 665938 24866 666174
rect 25102 665938 25134 666174
rect 24514 665854 25134 665938
rect 24514 665618 24546 665854
rect 24782 665618 24866 665854
rect 25102 665618 25134 665854
rect 24514 626174 25134 665618
rect 24514 625938 24546 626174
rect 24782 625938 24866 626174
rect 25102 625938 25134 626174
rect 24514 625854 25134 625938
rect 24514 625618 24546 625854
rect 24782 625618 24866 625854
rect 25102 625618 25134 625854
rect 24514 586174 25134 625618
rect 24514 585938 24546 586174
rect 24782 585938 24866 586174
rect 25102 585938 25134 586174
rect 24514 585854 25134 585938
rect 24514 585618 24546 585854
rect 24782 585618 24866 585854
rect 25102 585618 25134 585854
rect 24514 546174 25134 585618
rect 24514 545938 24546 546174
rect 24782 545938 24866 546174
rect 25102 545938 25134 546174
rect 24514 545854 25134 545938
rect 24514 545618 24546 545854
rect 24782 545618 24866 545854
rect 25102 545618 25134 545854
rect 24514 506174 25134 545618
rect 24514 505938 24546 506174
rect 24782 505938 24866 506174
rect 25102 505938 25134 506174
rect 24514 505854 25134 505938
rect 24514 505618 24546 505854
rect 24782 505618 24866 505854
rect 25102 505618 25134 505854
rect 24514 466174 25134 505618
rect 24514 465938 24546 466174
rect 24782 465938 24866 466174
rect 25102 465938 25134 466174
rect 24514 465854 25134 465938
rect 24514 465618 24546 465854
rect 24782 465618 24866 465854
rect 25102 465618 25134 465854
rect 24514 426174 25134 465618
rect 24514 425938 24546 426174
rect 24782 425938 24866 426174
rect 25102 425938 25134 426174
rect 24514 425854 25134 425938
rect 24514 425618 24546 425854
rect 24782 425618 24866 425854
rect 25102 425618 25134 425854
rect 24514 386174 25134 425618
rect 24514 385938 24546 386174
rect 24782 385938 24866 386174
rect 25102 385938 25134 386174
rect 24514 385854 25134 385938
rect 24514 385618 24546 385854
rect 24782 385618 24866 385854
rect 25102 385618 25134 385854
rect 24514 346174 25134 385618
rect 24514 345938 24546 346174
rect 24782 345938 24866 346174
rect 25102 345938 25134 346174
rect 24514 345854 25134 345938
rect 24514 345618 24546 345854
rect 24782 345618 24866 345854
rect 25102 345618 25134 345854
rect 24514 306174 25134 345618
rect 24514 305938 24546 306174
rect 24782 305938 24866 306174
rect 25102 305938 25134 306174
rect 24514 305854 25134 305938
rect 24514 305618 24546 305854
rect 24782 305618 24866 305854
rect 25102 305618 25134 305854
rect 24514 266174 25134 305618
rect 24514 265938 24546 266174
rect 24782 265938 24866 266174
rect 25102 265938 25134 266174
rect 24514 265854 25134 265938
rect 24514 265618 24546 265854
rect 24782 265618 24866 265854
rect 25102 265618 25134 265854
rect 24514 226174 25134 265618
rect 24514 225938 24546 226174
rect 24782 225938 24866 226174
rect 25102 225938 25134 226174
rect 24514 225854 25134 225938
rect 24514 225618 24546 225854
rect 24782 225618 24866 225854
rect 25102 225618 25134 225854
rect 24514 186174 25134 225618
rect 24514 185938 24546 186174
rect 24782 185938 24866 186174
rect 25102 185938 25134 186174
rect 24514 185854 25134 185938
rect 24514 185618 24546 185854
rect 24782 185618 24866 185854
rect 25102 185618 25134 185854
rect 24514 146174 25134 185618
rect 24514 145938 24546 146174
rect 24782 145938 24866 146174
rect 25102 145938 25134 146174
rect 24514 145854 25134 145938
rect 24514 145618 24546 145854
rect 24782 145618 24866 145854
rect 25102 145618 25134 145854
rect 24514 106174 25134 145618
rect 24514 105938 24546 106174
rect 24782 105938 24866 106174
rect 25102 105938 25134 106174
rect 24514 105854 25134 105938
rect 24514 105618 24546 105854
rect 24782 105618 24866 105854
rect 25102 105618 25134 105854
rect 24514 66174 25134 105618
rect 24514 65938 24546 66174
rect 24782 65938 24866 66174
rect 25102 65938 25134 66174
rect 24514 65854 25134 65938
rect 24514 65618 24546 65854
rect 24782 65618 24866 65854
rect 25102 65618 25134 65854
rect 24514 26174 25134 65618
rect 24514 25938 24546 26174
rect 24782 25938 24866 26174
rect 25102 25938 25134 26174
rect 24514 25854 25134 25938
rect 24514 25618 24546 25854
rect 24782 25618 24866 25854
rect 25102 25618 25134 25854
rect 24514 -3226 25134 25618
rect 24514 -3462 24546 -3226
rect 24782 -3462 24866 -3226
rect 25102 -3462 25134 -3226
rect 24514 -3546 25134 -3462
rect 24514 -3782 24546 -3546
rect 24782 -3782 24866 -3546
rect 25102 -3782 25134 -3546
rect 24514 -3814 25134 -3782
rect 28234 669894 28854 709082
rect 28234 669658 28266 669894
rect 28502 669658 28586 669894
rect 28822 669658 28854 669894
rect 28234 669574 28854 669658
rect 28234 669338 28266 669574
rect 28502 669338 28586 669574
rect 28822 669338 28854 669574
rect 28234 629894 28854 669338
rect 28234 629658 28266 629894
rect 28502 629658 28586 629894
rect 28822 629658 28854 629894
rect 28234 629574 28854 629658
rect 28234 629338 28266 629574
rect 28502 629338 28586 629574
rect 28822 629338 28854 629574
rect 28234 589894 28854 629338
rect 28234 589658 28266 589894
rect 28502 589658 28586 589894
rect 28822 589658 28854 589894
rect 28234 589574 28854 589658
rect 28234 589338 28266 589574
rect 28502 589338 28586 589574
rect 28822 589338 28854 589574
rect 28234 549894 28854 589338
rect 28234 549658 28266 549894
rect 28502 549658 28586 549894
rect 28822 549658 28854 549894
rect 28234 549574 28854 549658
rect 28234 549338 28266 549574
rect 28502 549338 28586 549574
rect 28822 549338 28854 549574
rect 28234 509894 28854 549338
rect 28234 509658 28266 509894
rect 28502 509658 28586 509894
rect 28822 509658 28854 509894
rect 28234 509574 28854 509658
rect 28234 509338 28266 509574
rect 28502 509338 28586 509574
rect 28822 509338 28854 509574
rect 28234 469894 28854 509338
rect 28234 469658 28266 469894
rect 28502 469658 28586 469894
rect 28822 469658 28854 469894
rect 28234 469574 28854 469658
rect 28234 469338 28266 469574
rect 28502 469338 28586 469574
rect 28822 469338 28854 469574
rect 28234 429894 28854 469338
rect 28234 429658 28266 429894
rect 28502 429658 28586 429894
rect 28822 429658 28854 429894
rect 28234 429574 28854 429658
rect 28234 429338 28266 429574
rect 28502 429338 28586 429574
rect 28822 429338 28854 429574
rect 28234 389894 28854 429338
rect 28234 389658 28266 389894
rect 28502 389658 28586 389894
rect 28822 389658 28854 389894
rect 28234 389574 28854 389658
rect 28234 389338 28266 389574
rect 28502 389338 28586 389574
rect 28822 389338 28854 389574
rect 28234 349894 28854 389338
rect 28234 349658 28266 349894
rect 28502 349658 28586 349894
rect 28822 349658 28854 349894
rect 28234 349574 28854 349658
rect 28234 349338 28266 349574
rect 28502 349338 28586 349574
rect 28822 349338 28854 349574
rect 28234 309894 28854 349338
rect 28234 309658 28266 309894
rect 28502 309658 28586 309894
rect 28822 309658 28854 309894
rect 28234 309574 28854 309658
rect 28234 309338 28266 309574
rect 28502 309338 28586 309574
rect 28822 309338 28854 309574
rect 28234 269894 28854 309338
rect 28234 269658 28266 269894
rect 28502 269658 28586 269894
rect 28822 269658 28854 269894
rect 28234 269574 28854 269658
rect 28234 269338 28266 269574
rect 28502 269338 28586 269574
rect 28822 269338 28854 269574
rect 28234 229894 28854 269338
rect 28234 229658 28266 229894
rect 28502 229658 28586 229894
rect 28822 229658 28854 229894
rect 28234 229574 28854 229658
rect 28234 229338 28266 229574
rect 28502 229338 28586 229574
rect 28822 229338 28854 229574
rect 28234 189894 28854 229338
rect 28234 189658 28266 189894
rect 28502 189658 28586 189894
rect 28822 189658 28854 189894
rect 28234 189574 28854 189658
rect 28234 189338 28266 189574
rect 28502 189338 28586 189574
rect 28822 189338 28854 189574
rect 28234 149894 28854 189338
rect 28234 149658 28266 149894
rect 28502 149658 28586 149894
rect 28822 149658 28854 149894
rect 28234 149574 28854 149658
rect 28234 149338 28266 149574
rect 28502 149338 28586 149574
rect 28822 149338 28854 149574
rect 28234 109894 28854 149338
rect 28234 109658 28266 109894
rect 28502 109658 28586 109894
rect 28822 109658 28854 109894
rect 28234 109574 28854 109658
rect 28234 109338 28266 109574
rect 28502 109338 28586 109574
rect 28822 109338 28854 109574
rect 28234 69894 28854 109338
rect 28234 69658 28266 69894
rect 28502 69658 28586 69894
rect 28822 69658 28854 69894
rect 28234 69574 28854 69658
rect 28234 69338 28266 69574
rect 28502 69338 28586 69574
rect 28822 69338 28854 69574
rect 28234 29894 28854 69338
rect 28234 29658 28266 29894
rect 28502 29658 28586 29894
rect 28822 29658 28854 29894
rect 28234 29574 28854 29658
rect 28234 29338 28266 29574
rect 28502 29338 28586 29574
rect 28822 29338 28854 29574
rect 28234 -5146 28854 29338
rect 28234 -5382 28266 -5146
rect 28502 -5382 28586 -5146
rect 28822 -5382 28854 -5146
rect 28234 -5466 28854 -5382
rect 28234 -5702 28266 -5466
rect 28502 -5702 28586 -5466
rect 28822 -5702 28854 -5466
rect 28234 -5734 28854 -5702
rect 31954 673614 32574 711002
rect 51954 710598 52574 711590
rect 51954 710362 51986 710598
rect 52222 710362 52306 710598
rect 52542 710362 52574 710598
rect 51954 710278 52574 710362
rect 51954 710042 51986 710278
rect 52222 710042 52306 710278
rect 52542 710042 52574 710278
rect 48234 708678 48854 709670
rect 48234 708442 48266 708678
rect 48502 708442 48586 708678
rect 48822 708442 48854 708678
rect 48234 708358 48854 708442
rect 48234 708122 48266 708358
rect 48502 708122 48586 708358
rect 48822 708122 48854 708358
rect 44514 706758 45134 707750
rect 44514 706522 44546 706758
rect 44782 706522 44866 706758
rect 45102 706522 45134 706758
rect 44514 706438 45134 706522
rect 44514 706202 44546 706438
rect 44782 706202 44866 706438
rect 45102 706202 45134 706438
rect 31954 673378 31986 673614
rect 32222 673378 32306 673614
rect 32542 673378 32574 673614
rect 31954 673294 32574 673378
rect 31954 673058 31986 673294
rect 32222 673058 32306 673294
rect 32542 673058 32574 673294
rect 31954 633614 32574 673058
rect 31954 633378 31986 633614
rect 32222 633378 32306 633614
rect 32542 633378 32574 633614
rect 31954 633294 32574 633378
rect 31954 633058 31986 633294
rect 32222 633058 32306 633294
rect 32542 633058 32574 633294
rect 31954 593614 32574 633058
rect 31954 593378 31986 593614
rect 32222 593378 32306 593614
rect 32542 593378 32574 593614
rect 31954 593294 32574 593378
rect 31954 593058 31986 593294
rect 32222 593058 32306 593294
rect 32542 593058 32574 593294
rect 31954 553614 32574 593058
rect 31954 553378 31986 553614
rect 32222 553378 32306 553614
rect 32542 553378 32574 553614
rect 31954 553294 32574 553378
rect 31954 553058 31986 553294
rect 32222 553058 32306 553294
rect 32542 553058 32574 553294
rect 31954 513614 32574 553058
rect 31954 513378 31986 513614
rect 32222 513378 32306 513614
rect 32542 513378 32574 513614
rect 31954 513294 32574 513378
rect 31954 513058 31986 513294
rect 32222 513058 32306 513294
rect 32542 513058 32574 513294
rect 31954 473614 32574 513058
rect 31954 473378 31986 473614
rect 32222 473378 32306 473614
rect 32542 473378 32574 473614
rect 31954 473294 32574 473378
rect 31954 473058 31986 473294
rect 32222 473058 32306 473294
rect 32542 473058 32574 473294
rect 31954 433614 32574 473058
rect 31954 433378 31986 433614
rect 32222 433378 32306 433614
rect 32542 433378 32574 433614
rect 31954 433294 32574 433378
rect 31954 433058 31986 433294
rect 32222 433058 32306 433294
rect 32542 433058 32574 433294
rect 31954 393614 32574 433058
rect 31954 393378 31986 393614
rect 32222 393378 32306 393614
rect 32542 393378 32574 393614
rect 31954 393294 32574 393378
rect 31954 393058 31986 393294
rect 32222 393058 32306 393294
rect 32542 393058 32574 393294
rect 31954 353614 32574 393058
rect 31954 353378 31986 353614
rect 32222 353378 32306 353614
rect 32542 353378 32574 353614
rect 31954 353294 32574 353378
rect 31954 353058 31986 353294
rect 32222 353058 32306 353294
rect 32542 353058 32574 353294
rect 31954 313614 32574 353058
rect 31954 313378 31986 313614
rect 32222 313378 32306 313614
rect 32542 313378 32574 313614
rect 31954 313294 32574 313378
rect 31954 313058 31986 313294
rect 32222 313058 32306 313294
rect 32542 313058 32574 313294
rect 31954 273614 32574 313058
rect 31954 273378 31986 273614
rect 32222 273378 32306 273614
rect 32542 273378 32574 273614
rect 31954 273294 32574 273378
rect 31954 273058 31986 273294
rect 32222 273058 32306 273294
rect 32542 273058 32574 273294
rect 31954 233614 32574 273058
rect 31954 233378 31986 233614
rect 32222 233378 32306 233614
rect 32542 233378 32574 233614
rect 31954 233294 32574 233378
rect 31954 233058 31986 233294
rect 32222 233058 32306 233294
rect 32542 233058 32574 233294
rect 31954 193614 32574 233058
rect 31954 193378 31986 193614
rect 32222 193378 32306 193614
rect 32542 193378 32574 193614
rect 31954 193294 32574 193378
rect 31954 193058 31986 193294
rect 32222 193058 32306 193294
rect 32542 193058 32574 193294
rect 31954 153614 32574 193058
rect 31954 153378 31986 153614
rect 32222 153378 32306 153614
rect 32542 153378 32574 153614
rect 31954 153294 32574 153378
rect 31954 153058 31986 153294
rect 32222 153058 32306 153294
rect 32542 153058 32574 153294
rect 31954 113614 32574 153058
rect 31954 113378 31986 113614
rect 32222 113378 32306 113614
rect 32542 113378 32574 113614
rect 31954 113294 32574 113378
rect 31954 113058 31986 113294
rect 32222 113058 32306 113294
rect 32542 113058 32574 113294
rect 31954 73614 32574 113058
rect 31954 73378 31986 73614
rect 32222 73378 32306 73614
rect 32542 73378 32574 73614
rect 31954 73294 32574 73378
rect 31954 73058 31986 73294
rect 32222 73058 32306 73294
rect 32542 73058 32574 73294
rect 31954 33614 32574 73058
rect 31954 33378 31986 33614
rect 32222 33378 32306 33614
rect 32542 33378 32574 33614
rect 31954 33294 32574 33378
rect 31954 33058 31986 33294
rect 32222 33058 32306 33294
rect 32542 33058 32574 33294
rect 11954 -6342 11986 -6106
rect 12222 -6342 12306 -6106
rect 12542 -6342 12574 -6106
rect 11954 -6426 12574 -6342
rect 11954 -6662 11986 -6426
rect 12222 -6662 12306 -6426
rect 12542 -6662 12574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 11954 -7654 12574 -6662
rect 31954 -7066 32574 33058
rect 40794 704838 41414 705830
rect 40794 704602 40826 704838
rect 41062 704602 41146 704838
rect 41382 704602 41414 704838
rect 40794 704518 41414 704602
rect 40794 704282 40826 704518
rect 41062 704282 41146 704518
rect 41382 704282 41414 704518
rect 40794 682454 41414 704282
rect 40794 682218 40826 682454
rect 41062 682218 41146 682454
rect 41382 682218 41414 682454
rect 40794 682134 41414 682218
rect 40794 681898 40826 682134
rect 41062 681898 41146 682134
rect 41382 681898 41414 682134
rect 40794 642454 41414 681898
rect 40794 642218 40826 642454
rect 41062 642218 41146 642454
rect 41382 642218 41414 642454
rect 40794 642134 41414 642218
rect 40794 641898 40826 642134
rect 41062 641898 41146 642134
rect 41382 641898 41414 642134
rect 40794 602454 41414 641898
rect 40794 602218 40826 602454
rect 41062 602218 41146 602454
rect 41382 602218 41414 602454
rect 40794 602134 41414 602218
rect 40794 601898 40826 602134
rect 41062 601898 41146 602134
rect 41382 601898 41414 602134
rect 40794 562454 41414 601898
rect 40794 562218 40826 562454
rect 41062 562218 41146 562454
rect 41382 562218 41414 562454
rect 40794 562134 41414 562218
rect 40794 561898 40826 562134
rect 41062 561898 41146 562134
rect 41382 561898 41414 562134
rect 40794 522454 41414 561898
rect 40794 522218 40826 522454
rect 41062 522218 41146 522454
rect 41382 522218 41414 522454
rect 40794 522134 41414 522218
rect 40794 521898 40826 522134
rect 41062 521898 41146 522134
rect 41382 521898 41414 522134
rect 40794 482454 41414 521898
rect 40794 482218 40826 482454
rect 41062 482218 41146 482454
rect 41382 482218 41414 482454
rect 40794 482134 41414 482218
rect 40794 481898 40826 482134
rect 41062 481898 41146 482134
rect 41382 481898 41414 482134
rect 40794 442454 41414 481898
rect 40794 442218 40826 442454
rect 41062 442218 41146 442454
rect 41382 442218 41414 442454
rect 40794 442134 41414 442218
rect 40794 441898 40826 442134
rect 41062 441898 41146 442134
rect 41382 441898 41414 442134
rect 40794 402454 41414 441898
rect 40794 402218 40826 402454
rect 41062 402218 41146 402454
rect 41382 402218 41414 402454
rect 40794 402134 41414 402218
rect 40794 401898 40826 402134
rect 41062 401898 41146 402134
rect 41382 401898 41414 402134
rect 40794 362454 41414 401898
rect 40794 362218 40826 362454
rect 41062 362218 41146 362454
rect 41382 362218 41414 362454
rect 40794 362134 41414 362218
rect 40794 361898 40826 362134
rect 41062 361898 41146 362134
rect 41382 361898 41414 362134
rect 40794 322454 41414 361898
rect 40794 322218 40826 322454
rect 41062 322218 41146 322454
rect 41382 322218 41414 322454
rect 40794 322134 41414 322218
rect 40794 321898 40826 322134
rect 41062 321898 41146 322134
rect 41382 321898 41414 322134
rect 40794 282454 41414 321898
rect 40794 282218 40826 282454
rect 41062 282218 41146 282454
rect 41382 282218 41414 282454
rect 40794 282134 41414 282218
rect 40794 281898 40826 282134
rect 41062 281898 41146 282134
rect 41382 281898 41414 282134
rect 40794 242454 41414 281898
rect 40794 242218 40826 242454
rect 41062 242218 41146 242454
rect 41382 242218 41414 242454
rect 40794 242134 41414 242218
rect 40794 241898 40826 242134
rect 41062 241898 41146 242134
rect 41382 241898 41414 242134
rect 40794 202454 41414 241898
rect 40794 202218 40826 202454
rect 41062 202218 41146 202454
rect 41382 202218 41414 202454
rect 40794 202134 41414 202218
rect 40794 201898 40826 202134
rect 41062 201898 41146 202134
rect 41382 201898 41414 202134
rect 40794 162454 41414 201898
rect 40794 162218 40826 162454
rect 41062 162218 41146 162454
rect 41382 162218 41414 162454
rect 40794 162134 41414 162218
rect 40794 161898 40826 162134
rect 41062 161898 41146 162134
rect 41382 161898 41414 162134
rect 40794 122454 41414 161898
rect 40794 122218 40826 122454
rect 41062 122218 41146 122454
rect 41382 122218 41414 122454
rect 40794 122134 41414 122218
rect 40794 121898 40826 122134
rect 41062 121898 41146 122134
rect 41382 121898 41414 122134
rect 40794 82454 41414 121898
rect 40794 82218 40826 82454
rect 41062 82218 41146 82454
rect 41382 82218 41414 82454
rect 40794 82134 41414 82218
rect 40794 81898 40826 82134
rect 41062 81898 41146 82134
rect 41382 81898 41414 82134
rect 40794 42454 41414 81898
rect 40794 42218 40826 42454
rect 41062 42218 41146 42454
rect 41382 42218 41414 42454
rect 40794 42134 41414 42218
rect 40794 41898 40826 42134
rect 41062 41898 41146 42134
rect 41382 41898 41414 42134
rect 40794 2454 41414 41898
rect 40794 2218 40826 2454
rect 41062 2218 41146 2454
rect 41382 2218 41414 2454
rect 40794 2134 41414 2218
rect 40794 1898 40826 2134
rect 41062 1898 41146 2134
rect 41382 1898 41414 2134
rect 40794 -346 41414 1898
rect 40794 -582 40826 -346
rect 41062 -582 41146 -346
rect 41382 -582 41414 -346
rect 40794 -666 41414 -582
rect 40794 -902 40826 -666
rect 41062 -902 41146 -666
rect 41382 -902 41414 -666
rect 40794 -1894 41414 -902
rect 44514 686174 45134 706202
rect 44514 685938 44546 686174
rect 44782 685938 44866 686174
rect 45102 685938 45134 686174
rect 44514 685854 45134 685938
rect 44514 685618 44546 685854
rect 44782 685618 44866 685854
rect 45102 685618 45134 685854
rect 44514 646174 45134 685618
rect 44514 645938 44546 646174
rect 44782 645938 44866 646174
rect 45102 645938 45134 646174
rect 44514 645854 45134 645938
rect 44514 645618 44546 645854
rect 44782 645618 44866 645854
rect 45102 645618 45134 645854
rect 44514 606174 45134 645618
rect 44514 605938 44546 606174
rect 44782 605938 44866 606174
rect 45102 605938 45134 606174
rect 44514 605854 45134 605938
rect 44514 605618 44546 605854
rect 44782 605618 44866 605854
rect 45102 605618 45134 605854
rect 44514 566174 45134 605618
rect 44514 565938 44546 566174
rect 44782 565938 44866 566174
rect 45102 565938 45134 566174
rect 44514 565854 45134 565938
rect 44514 565618 44546 565854
rect 44782 565618 44866 565854
rect 45102 565618 45134 565854
rect 44514 526174 45134 565618
rect 44514 525938 44546 526174
rect 44782 525938 44866 526174
rect 45102 525938 45134 526174
rect 44514 525854 45134 525938
rect 44514 525618 44546 525854
rect 44782 525618 44866 525854
rect 45102 525618 45134 525854
rect 44514 486174 45134 525618
rect 44514 485938 44546 486174
rect 44782 485938 44866 486174
rect 45102 485938 45134 486174
rect 44514 485854 45134 485938
rect 44514 485618 44546 485854
rect 44782 485618 44866 485854
rect 45102 485618 45134 485854
rect 44514 446174 45134 485618
rect 44514 445938 44546 446174
rect 44782 445938 44866 446174
rect 45102 445938 45134 446174
rect 44514 445854 45134 445938
rect 44514 445618 44546 445854
rect 44782 445618 44866 445854
rect 45102 445618 45134 445854
rect 44514 406174 45134 445618
rect 44514 405938 44546 406174
rect 44782 405938 44866 406174
rect 45102 405938 45134 406174
rect 44514 405854 45134 405938
rect 44514 405618 44546 405854
rect 44782 405618 44866 405854
rect 45102 405618 45134 405854
rect 44514 366174 45134 405618
rect 44514 365938 44546 366174
rect 44782 365938 44866 366174
rect 45102 365938 45134 366174
rect 44514 365854 45134 365938
rect 44514 365618 44546 365854
rect 44782 365618 44866 365854
rect 45102 365618 45134 365854
rect 44514 326174 45134 365618
rect 44514 325938 44546 326174
rect 44782 325938 44866 326174
rect 45102 325938 45134 326174
rect 44514 325854 45134 325938
rect 44514 325618 44546 325854
rect 44782 325618 44866 325854
rect 45102 325618 45134 325854
rect 44514 286174 45134 325618
rect 44514 285938 44546 286174
rect 44782 285938 44866 286174
rect 45102 285938 45134 286174
rect 44514 285854 45134 285938
rect 44514 285618 44546 285854
rect 44782 285618 44866 285854
rect 45102 285618 45134 285854
rect 44514 246174 45134 285618
rect 44514 245938 44546 246174
rect 44782 245938 44866 246174
rect 45102 245938 45134 246174
rect 44514 245854 45134 245938
rect 44514 245618 44546 245854
rect 44782 245618 44866 245854
rect 45102 245618 45134 245854
rect 44514 206174 45134 245618
rect 44514 205938 44546 206174
rect 44782 205938 44866 206174
rect 45102 205938 45134 206174
rect 44514 205854 45134 205938
rect 44514 205618 44546 205854
rect 44782 205618 44866 205854
rect 45102 205618 45134 205854
rect 44514 166174 45134 205618
rect 44514 165938 44546 166174
rect 44782 165938 44866 166174
rect 45102 165938 45134 166174
rect 44514 165854 45134 165938
rect 44514 165618 44546 165854
rect 44782 165618 44866 165854
rect 45102 165618 45134 165854
rect 44514 126174 45134 165618
rect 44514 125938 44546 126174
rect 44782 125938 44866 126174
rect 45102 125938 45134 126174
rect 44514 125854 45134 125938
rect 44514 125618 44546 125854
rect 44782 125618 44866 125854
rect 45102 125618 45134 125854
rect 44514 86174 45134 125618
rect 44514 85938 44546 86174
rect 44782 85938 44866 86174
rect 45102 85938 45134 86174
rect 44514 85854 45134 85938
rect 44514 85618 44546 85854
rect 44782 85618 44866 85854
rect 45102 85618 45134 85854
rect 44514 46174 45134 85618
rect 44514 45938 44546 46174
rect 44782 45938 44866 46174
rect 45102 45938 45134 46174
rect 44514 45854 45134 45938
rect 44514 45618 44546 45854
rect 44782 45618 44866 45854
rect 45102 45618 45134 45854
rect 44514 6174 45134 45618
rect 44514 5938 44546 6174
rect 44782 5938 44866 6174
rect 45102 5938 45134 6174
rect 44514 5854 45134 5938
rect 44514 5618 44546 5854
rect 44782 5618 44866 5854
rect 45102 5618 45134 5854
rect 44514 -2266 45134 5618
rect 44514 -2502 44546 -2266
rect 44782 -2502 44866 -2266
rect 45102 -2502 45134 -2266
rect 44514 -2586 45134 -2502
rect 44514 -2822 44546 -2586
rect 44782 -2822 44866 -2586
rect 45102 -2822 45134 -2586
rect 44514 -3814 45134 -2822
rect 48234 689894 48854 708122
rect 48234 689658 48266 689894
rect 48502 689658 48586 689894
rect 48822 689658 48854 689894
rect 48234 689574 48854 689658
rect 48234 689338 48266 689574
rect 48502 689338 48586 689574
rect 48822 689338 48854 689574
rect 48234 649894 48854 689338
rect 48234 649658 48266 649894
rect 48502 649658 48586 649894
rect 48822 649658 48854 649894
rect 48234 649574 48854 649658
rect 48234 649338 48266 649574
rect 48502 649338 48586 649574
rect 48822 649338 48854 649574
rect 48234 609894 48854 649338
rect 48234 609658 48266 609894
rect 48502 609658 48586 609894
rect 48822 609658 48854 609894
rect 48234 609574 48854 609658
rect 48234 609338 48266 609574
rect 48502 609338 48586 609574
rect 48822 609338 48854 609574
rect 48234 569894 48854 609338
rect 48234 569658 48266 569894
rect 48502 569658 48586 569894
rect 48822 569658 48854 569894
rect 48234 569574 48854 569658
rect 48234 569338 48266 569574
rect 48502 569338 48586 569574
rect 48822 569338 48854 569574
rect 48234 529894 48854 569338
rect 48234 529658 48266 529894
rect 48502 529658 48586 529894
rect 48822 529658 48854 529894
rect 48234 529574 48854 529658
rect 48234 529338 48266 529574
rect 48502 529338 48586 529574
rect 48822 529338 48854 529574
rect 48234 489894 48854 529338
rect 48234 489658 48266 489894
rect 48502 489658 48586 489894
rect 48822 489658 48854 489894
rect 48234 489574 48854 489658
rect 48234 489338 48266 489574
rect 48502 489338 48586 489574
rect 48822 489338 48854 489574
rect 48234 449894 48854 489338
rect 48234 449658 48266 449894
rect 48502 449658 48586 449894
rect 48822 449658 48854 449894
rect 48234 449574 48854 449658
rect 48234 449338 48266 449574
rect 48502 449338 48586 449574
rect 48822 449338 48854 449574
rect 48234 409894 48854 449338
rect 48234 409658 48266 409894
rect 48502 409658 48586 409894
rect 48822 409658 48854 409894
rect 48234 409574 48854 409658
rect 48234 409338 48266 409574
rect 48502 409338 48586 409574
rect 48822 409338 48854 409574
rect 48234 369894 48854 409338
rect 48234 369658 48266 369894
rect 48502 369658 48586 369894
rect 48822 369658 48854 369894
rect 48234 369574 48854 369658
rect 48234 369338 48266 369574
rect 48502 369338 48586 369574
rect 48822 369338 48854 369574
rect 48234 329894 48854 369338
rect 48234 329658 48266 329894
rect 48502 329658 48586 329894
rect 48822 329658 48854 329894
rect 48234 329574 48854 329658
rect 48234 329338 48266 329574
rect 48502 329338 48586 329574
rect 48822 329338 48854 329574
rect 48234 289894 48854 329338
rect 48234 289658 48266 289894
rect 48502 289658 48586 289894
rect 48822 289658 48854 289894
rect 48234 289574 48854 289658
rect 48234 289338 48266 289574
rect 48502 289338 48586 289574
rect 48822 289338 48854 289574
rect 48234 249894 48854 289338
rect 48234 249658 48266 249894
rect 48502 249658 48586 249894
rect 48822 249658 48854 249894
rect 48234 249574 48854 249658
rect 48234 249338 48266 249574
rect 48502 249338 48586 249574
rect 48822 249338 48854 249574
rect 48234 209894 48854 249338
rect 48234 209658 48266 209894
rect 48502 209658 48586 209894
rect 48822 209658 48854 209894
rect 48234 209574 48854 209658
rect 48234 209338 48266 209574
rect 48502 209338 48586 209574
rect 48822 209338 48854 209574
rect 48234 169894 48854 209338
rect 48234 169658 48266 169894
rect 48502 169658 48586 169894
rect 48822 169658 48854 169894
rect 48234 169574 48854 169658
rect 48234 169338 48266 169574
rect 48502 169338 48586 169574
rect 48822 169338 48854 169574
rect 48234 129894 48854 169338
rect 48234 129658 48266 129894
rect 48502 129658 48586 129894
rect 48822 129658 48854 129894
rect 48234 129574 48854 129658
rect 48234 129338 48266 129574
rect 48502 129338 48586 129574
rect 48822 129338 48854 129574
rect 48234 89894 48854 129338
rect 48234 89658 48266 89894
rect 48502 89658 48586 89894
rect 48822 89658 48854 89894
rect 48234 89574 48854 89658
rect 48234 89338 48266 89574
rect 48502 89338 48586 89574
rect 48822 89338 48854 89574
rect 48234 49894 48854 89338
rect 48234 49658 48266 49894
rect 48502 49658 48586 49894
rect 48822 49658 48854 49894
rect 48234 49574 48854 49658
rect 48234 49338 48266 49574
rect 48502 49338 48586 49574
rect 48822 49338 48854 49574
rect 48234 9894 48854 49338
rect 48234 9658 48266 9894
rect 48502 9658 48586 9894
rect 48822 9658 48854 9894
rect 48234 9574 48854 9658
rect 48234 9338 48266 9574
rect 48502 9338 48586 9574
rect 48822 9338 48854 9574
rect 48234 -4186 48854 9338
rect 48234 -4422 48266 -4186
rect 48502 -4422 48586 -4186
rect 48822 -4422 48854 -4186
rect 48234 -4506 48854 -4422
rect 48234 -4742 48266 -4506
rect 48502 -4742 48586 -4506
rect 48822 -4742 48854 -4506
rect 48234 -5734 48854 -4742
rect 51954 693614 52574 710042
rect 71954 711558 72574 711590
rect 71954 711322 71986 711558
rect 72222 711322 72306 711558
rect 72542 711322 72574 711558
rect 71954 711238 72574 711322
rect 71954 711002 71986 711238
rect 72222 711002 72306 711238
rect 72542 711002 72574 711238
rect 68234 709638 68854 709670
rect 68234 709402 68266 709638
rect 68502 709402 68586 709638
rect 68822 709402 68854 709638
rect 68234 709318 68854 709402
rect 68234 709082 68266 709318
rect 68502 709082 68586 709318
rect 68822 709082 68854 709318
rect 64514 707718 65134 707750
rect 64514 707482 64546 707718
rect 64782 707482 64866 707718
rect 65102 707482 65134 707718
rect 64514 707398 65134 707482
rect 64514 707162 64546 707398
rect 64782 707162 64866 707398
rect 65102 707162 65134 707398
rect 51954 693378 51986 693614
rect 52222 693378 52306 693614
rect 52542 693378 52574 693614
rect 51954 693294 52574 693378
rect 51954 693058 51986 693294
rect 52222 693058 52306 693294
rect 52542 693058 52574 693294
rect 51954 653614 52574 693058
rect 51954 653378 51986 653614
rect 52222 653378 52306 653614
rect 52542 653378 52574 653614
rect 51954 653294 52574 653378
rect 51954 653058 51986 653294
rect 52222 653058 52306 653294
rect 52542 653058 52574 653294
rect 51954 613614 52574 653058
rect 51954 613378 51986 613614
rect 52222 613378 52306 613614
rect 52542 613378 52574 613614
rect 51954 613294 52574 613378
rect 51954 613058 51986 613294
rect 52222 613058 52306 613294
rect 52542 613058 52574 613294
rect 51954 573614 52574 613058
rect 51954 573378 51986 573614
rect 52222 573378 52306 573614
rect 52542 573378 52574 573614
rect 51954 573294 52574 573378
rect 51954 573058 51986 573294
rect 52222 573058 52306 573294
rect 52542 573058 52574 573294
rect 51954 533614 52574 573058
rect 51954 533378 51986 533614
rect 52222 533378 52306 533614
rect 52542 533378 52574 533614
rect 51954 533294 52574 533378
rect 51954 533058 51986 533294
rect 52222 533058 52306 533294
rect 52542 533058 52574 533294
rect 51954 493614 52574 533058
rect 51954 493378 51986 493614
rect 52222 493378 52306 493614
rect 52542 493378 52574 493614
rect 51954 493294 52574 493378
rect 51954 493058 51986 493294
rect 52222 493058 52306 493294
rect 52542 493058 52574 493294
rect 51954 453614 52574 493058
rect 51954 453378 51986 453614
rect 52222 453378 52306 453614
rect 52542 453378 52574 453614
rect 51954 453294 52574 453378
rect 51954 453058 51986 453294
rect 52222 453058 52306 453294
rect 52542 453058 52574 453294
rect 51954 413614 52574 453058
rect 51954 413378 51986 413614
rect 52222 413378 52306 413614
rect 52542 413378 52574 413614
rect 51954 413294 52574 413378
rect 51954 413058 51986 413294
rect 52222 413058 52306 413294
rect 52542 413058 52574 413294
rect 51954 373614 52574 413058
rect 51954 373378 51986 373614
rect 52222 373378 52306 373614
rect 52542 373378 52574 373614
rect 51954 373294 52574 373378
rect 51954 373058 51986 373294
rect 52222 373058 52306 373294
rect 52542 373058 52574 373294
rect 51954 333614 52574 373058
rect 51954 333378 51986 333614
rect 52222 333378 52306 333614
rect 52542 333378 52574 333614
rect 51954 333294 52574 333378
rect 51954 333058 51986 333294
rect 52222 333058 52306 333294
rect 52542 333058 52574 333294
rect 51954 293614 52574 333058
rect 51954 293378 51986 293614
rect 52222 293378 52306 293614
rect 52542 293378 52574 293614
rect 51954 293294 52574 293378
rect 51954 293058 51986 293294
rect 52222 293058 52306 293294
rect 52542 293058 52574 293294
rect 51954 253614 52574 293058
rect 51954 253378 51986 253614
rect 52222 253378 52306 253614
rect 52542 253378 52574 253614
rect 51954 253294 52574 253378
rect 51954 253058 51986 253294
rect 52222 253058 52306 253294
rect 52542 253058 52574 253294
rect 51954 213614 52574 253058
rect 51954 213378 51986 213614
rect 52222 213378 52306 213614
rect 52542 213378 52574 213614
rect 51954 213294 52574 213378
rect 51954 213058 51986 213294
rect 52222 213058 52306 213294
rect 52542 213058 52574 213294
rect 51954 173614 52574 213058
rect 51954 173378 51986 173614
rect 52222 173378 52306 173614
rect 52542 173378 52574 173614
rect 51954 173294 52574 173378
rect 51954 173058 51986 173294
rect 52222 173058 52306 173294
rect 52542 173058 52574 173294
rect 51954 133614 52574 173058
rect 51954 133378 51986 133614
rect 52222 133378 52306 133614
rect 52542 133378 52574 133614
rect 51954 133294 52574 133378
rect 51954 133058 51986 133294
rect 52222 133058 52306 133294
rect 52542 133058 52574 133294
rect 51954 93614 52574 133058
rect 51954 93378 51986 93614
rect 52222 93378 52306 93614
rect 52542 93378 52574 93614
rect 51954 93294 52574 93378
rect 51954 93058 51986 93294
rect 52222 93058 52306 93294
rect 52542 93058 52574 93294
rect 51954 53614 52574 93058
rect 51954 53378 51986 53614
rect 52222 53378 52306 53614
rect 52542 53378 52574 53614
rect 51954 53294 52574 53378
rect 51954 53058 51986 53294
rect 52222 53058 52306 53294
rect 52542 53058 52574 53294
rect 51954 13614 52574 53058
rect 51954 13378 51986 13614
rect 52222 13378 52306 13614
rect 52542 13378 52574 13614
rect 51954 13294 52574 13378
rect 51954 13058 51986 13294
rect 52222 13058 52306 13294
rect 52542 13058 52574 13294
rect 31954 -7302 31986 -7066
rect 32222 -7302 32306 -7066
rect 32542 -7302 32574 -7066
rect 31954 -7386 32574 -7302
rect 31954 -7622 31986 -7386
rect 32222 -7622 32306 -7386
rect 32542 -7622 32574 -7386
rect 31954 -7654 32574 -7622
rect 51954 -6106 52574 13058
rect 60794 705798 61414 705830
rect 60794 705562 60826 705798
rect 61062 705562 61146 705798
rect 61382 705562 61414 705798
rect 60794 705478 61414 705562
rect 60794 705242 60826 705478
rect 61062 705242 61146 705478
rect 61382 705242 61414 705478
rect 60794 662454 61414 705242
rect 60794 662218 60826 662454
rect 61062 662218 61146 662454
rect 61382 662218 61414 662454
rect 60794 662134 61414 662218
rect 60794 661898 60826 662134
rect 61062 661898 61146 662134
rect 61382 661898 61414 662134
rect 60794 622454 61414 661898
rect 60794 622218 60826 622454
rect 61062 622218 61146 622454
rect 61382 622218 61414 622454
rect 60794 622134 61414 622218
rect 60794 621898 60826 622134
rect 61062 621898 61146 622134
rect 61382 621898 61414 622134
rect 60794 582454 61414 621898
rect 60794 582218 60826 582454
rect 61062 582218 61146 582454
rect 61382 582218 61414 582454
rect 60794 582134 61414 582218
rect 60794 581898 60826 582134
rect 61062 581898 61146 582134
rect 61382 581898 61414 582134
rect 60794 542454 61414 581898
rect 60794 542218 60826 542454
rect 61062 542218 61146 542454
rect 61382 542218 61414 542454
rect 60794 542134 61414 542218
rect 60794 541898 60826 542134
rect 61062 541898 61146 542134
rect 61382 541898 61414 542134
rect 60794 502454 61414 541898
rect 60794 502218 60826 502454
rect 61062 502218 61146 502454
rect 61382 502218 61414 502454
rect 60794 502134 61414 502218
rect 60794 501898 60826 502134
rect 61062 501898 61146 502134
rect 61382 501898 61414 502134
rect 60794 462454 61414 501898
rect 60794 462218 60826 462454
rect 61062 462218 61146 462454
rect 61382 462218 61414 462454
rect 60794 462134 61414 462218
rect 60794 461898 60826 462134
rect 61062 461898 61146 462134
rect 61382 461898 61414 462134
rect 60794 422454 61414 461898
rect 60794 422218 60826 422454
rect 61062 422218 61146 422454
rect 61382 422218 61414 422454
rect 60794 422134 61414 422218
rect 60794 421898 60826 422134
rect 61062 421898 61146 422134
rect 61382 421898 61414 422134
rect 60794 382454 61414 421898
rect 60794 382218 60826 382454
rect 61062 382218 61146 382454
rect 61382 382218 61414 382454
rect 60794 382134 61414 382218
rect 60794 381898 60826 382134
rect 61062 381898 61146 382134
rect 61382 381898 61414 382134
rect 60794 342454 61414 381898
rect 60794 342218 60826 342454
rect 61062 342218 61146 342454
rect 61382 342218 61414 342454
rect 60794 342134 61414 342218
rect 60794 341898 60826 342134
rect 61062 341898 61146 342134
rect 61382 341898 61414 342134
rect 60794 302454 61414 341898
rect 60794 302218 60826 302454
rect 61062 302218 61146 302454
rect 61382 302218 61414 302454
rect 60794 302134 61414 302218
rect 60794 301898 60826 302134
rect 61062 301898 61146 302134
rect 61382 301898 61414 302134
rect 60794 262454 61414 301898
rect 60794 262218 60826 262454
rect 61062 262218 61146 262454
rect 61382 262218 61414 262454
rect 60794 262134 61414 262218
rect 60794 261898 60826 262134
rect 61062 261898 61146 262134
rect 61382 261898 61414 262134
rect 60794 222454 61414 261898
rect 60794 222218 60826 222454
rect 61062 222218 61146 222454
rect 61382 222218 61414 222454
rect 60794 222134 61414 222218
rect 60794 221898 60826 222134
rect 61062 221898 61146 222134
rect 61382 221898 61414 222134
rect 60794 182454 61414 221898
rect 60794 182218 60826 182454
rect 61062 182218 61146 182454
rect 61382 182218 61414 182454
rect 60794 182134 61414 182218
rect 60794 181898 60826 182134
rect 61062 181898 61146 182134
rect 61382 181898 61414 182134
rect 60794 142454 61414 181898
rect 60794 142218 60826 142454
rect 61062 142218 61146 142454
rect 61382 142218 61414 142454
rect 60794 142134 61414 142218
rect 60794 141898 60826 142134
rect 61062 141898 61146 142134
rect 61382 141898 61414 142134
rect 60794 102454 61414 141898
rect 60794 102218 60826 102454
rect 61062 102218 61146 102454
rect 61382 102218 61414 102454
rect 60794 102134 61414 102218
rect 60794 101898 60826 102134
rect 61062 101898 61146 102134
rect 61382 101898 61414 102134
rect 60794 62454 61414 101898
rect 60794 62218 60826 62454
rect 61062 62218 61146 62454
rect 61382 62218 61414 62454
rect 60794 62134 61414 62218
rect 60794 61898 60826 62134
rect 61062 61898 61146 62134
rect 61382 61898 61414 62134
rect 60794 22454 61414 61898
rect 60794 22218 60826 22454
rect 61062 22218 61146 22454
rect 61382 22218 61414 22454
rect 60794 22134 61414 22218
rect 60794 21898 60826 22134
rect 61062 21898 61146 22134
rect 61382 21898 61414 22134
rect 60794 -1306 61414 21898
rect 60794 -1542 60826 -1306
rect 61062 -1542 61146 -1306
rect 61382 -1542 61414 -1306
rect 60794 -1626 61414 -1542
rect 60794 -1862 60826 -1626
rect 61062 -1862 61146 -1626
rect 61382 -1862 61414 -1626
rect 60794 -1894 61414 -1862
rect 64514 666174 65134 707162
rect 64514 665938 64546 666174
rect 64782 665938 64866 666174
rect 65102 665938 65134 666174
rect 64514 665854 65134 665938
rect 64514 665618 64546 665854
rect 64782 665618 64866 665854
rect 65102 665618 65134 665854
rect 64514 626174 65134 665618
rect 64514 625938 64546 626174
rect 64782 625938 64866 626174
rect 65102 625938 65134 626174
rect 64514 625854 65134 625938
rect 64514 625618 64546 625854
rect 64782 625618 64866 625854
rect 65102 625618 65134 625854
rect 64514 586174 65134 625618
rect 64514 585938 64546 586174
rect 64782 585938 64866 586174
rect 65102 585938 65134 586174
rect 64514 585854 65134 585938
rect 64514 585618 64546 585854
rect 64782 585618 64866 585854
rect 65102 585618 65134 585854
rect 64514 546174 65134 585618
rect 64514 545938 64546 546174
rect 64782 545938 64866 546174
rect 65102 545938 65134 546174
rect 64514 545854 65134 545938
rect 64514 545618 64546 545854
rect 64782 545618 64866 545854
rect 65102 545618 65134 545854
rect 64514 506174 65134 545618
rect 64514 505938 64546 506174
rect 64782 505938 64866 506174
rect 65102 505938 65134 506174
rect 64514 505854 65134 505938
rect 64514 505618 64546 505854
rect 64782 505618 64866 505854
rect 65102 505618 65134 505854
rect 64514 466174 65134 505618
rect 64514 465938 64546 466174
rect 64782 465938 64866 466174
rect 65102 465938 65134 466174
rect 64514 465854 65134 465938
rect 64514 465618 64546 465854
rect 64782 465618 64866 465854
rect 65102 465618 65134 465854
rect 64514 426174 65134 465618
rect 64514 425938 64546 426174
rect 64782 425938 64866 426174
rect 65102 425938 65134 426174
rect 64514 425854 65134 425938
rect 64514 425618 64546 425854
rect 64782 425618 64866 425854
rect 65102 425618 65134 425854
rect 64514 386174 65134 425618
rect 64514 385938 64546 386174
rect 64782 385938 64866 386174
rect 65102 385938 65134 386174
rect 64514 385854 65134 385938
rect 64514 385618 64546 385854
rect 64782 385618 64866 385854
rect 65102 385618 65134 385854
rect 64514 346174 65134 385618
rect 64514 345938 64546 346174
rect 64782 345938 64866 346174
rect 65102 345938 65134 346174
rect 64514 345854 65134 345938
rect 64514 345618 64546 345854
rect 64782 345618 64866 345854
rect 65102 345618 65134 345854
rect 64514 306174 65134 345618
rect 64514 305938 64546 306174
rect 64782 305938 64866 306174
rect 65102 305938 65134 306174
rect 64514 305854 65134 305938
rect 64514 305618 64546 305854
rect 64782 305618 64866 305854
rect 65102 305618 65134 305854
rect 64514 266174 65134 305618
rect 64514 265938 64546 266174
rect 64782 265938 64866 266174
rect 65102 265938 65134 266174
rect 64514 265854 65134 265938
rect 64514 265618 64546 265854
rect 64782 265618 64866 265854
rect 65102 265618 65134 265854
rect 64514 226174 65134 265618
rect 64514 225938 64546 226174
rect 64782 225938 64866 226174
rect 65102 225938 65134 226174
rect 64514 225854 65134 225938
rect 64514 225618 64546 225854
rect 64782 225618 64866 225854
rect 65102 225618 65134 225854
rect 64514 186174 65134 225618
rect 64514 185938 64546 186174
rect 64782 185938 64866 186174
rect 65102 185938 65134 186174
rect 64514 185854 65134 185938
rect 64514 185618 64546 185854
rect 64782 185618 64866 185854
rect 65102 185618 65134 185854
rect 64514 146174 65134 185618
rect 64514 145938 64546 146174
rect 64782 145938 64866 146174
rect 65102 145938 65134 146174
rect 64514 145854 65134 145938
rect 64514 145618 64546 145854
rect 64782 145618 64866 145854
rect 65102 145618 65134 145854
rect 64514 106174 65134 145618
rect 64514 105938 64546 106174
rect 64782 105938 64866 106174
rect 65102 105938 65134 106174
rect 64514 105854 65134 105938
rect 64514 105618 64546 105854
rect 64782 105618 64866 105854
rect 65102 105618 65134 105854
rect 64514 66174 65134 105618
rect 64514 65938 64546 66174
rect 64782 65938 64866 66174
rect 65102 65938 65134 66174
rect 64514 65854 65134 65938
rect 64514 65618 64546 65854
rect 64782 65618 64866 65854
rect 65102 65618 65134 65854
rect 64514 26174 65134 65618
rect 64514 25938 64546 26174
rect 64782 25938 64866 26174
rect 65102 25938 65134 26174
rect 64514 25854 65134 25938
rect 64514 25618 64546 25854
rect 64782 25618 64866 25854
rect 65102 25618 65134 25854
rect 64514 -3226 65134 25618
rect 64514 -3462 64546 -3226
rect 64782 -3462 64866 -3226
rect 65102 -3462 65134 -3226
rect 64514 -3546 65134 -3462
rect 64514 -3782 64546 -3546
rect 64782 -3782 64866 -3546
rect 65102 -3782 65134 -3546
rect 64514 -3814 65134 -3782
rect 68234 669894 68854 709082
rect 68234 669658 68266 669894
rect 68502 669658 68586 669894
rect 68822 669658 68854 669894
rect 68234 669574 68854 669658
rect 68234 669338 68266 669574
rect 68502 669338 68586 669574
rect 68822 669338 68854 669574
rect 68234 629894 68854 669338
rect 68234 629658 68266 629894
rect 68502 629658 68586 629894
rect 68822 629658 68854 629894
rect 68234 629574 68854 629658
rect 68234 629338 68266 629574
rect 68502 629338 68586 629574
rect 68822 629338 68854 629574
rect 68234 589894 68854 629338
rect 68234 589658 68266 589894
rect 68502 589658 68586 589894
rect 68822 589658 68854 589894
rect 68234 589574 68854 589658
rect 68234 589338 68266 589574
rect 68502 589338 68586 589574
rect 68822 589338 68854 589574
rect 68234 549894 68854 589338
rect 68234 549658 68266 549894
rect 68502 549658 68586 549894
rect 68822 549658 68854 549894
rect 68234 549574 68854 549658
rect 68234 549338 68266 549574
rect 68502 549338 68586 549574
rect 68822 549338 68854 549574
rect 68234 509894 68854 549338
rect 68234 509658 68266 509894
rect 68502 509658 68586 509894
rect 68822 509658 68854 509894
rect 68234 509574 68854 509658
rect 68234 509338 68266 509574
rect 68502 509338 68586 509574
rect 68822 509338 68854 509574
rect 68234 469894 68854 509338
rect 68234 469658 68266 469894
rect 68502 469658 68586 469894
rect 68822 469658 68854 469894
rect 68234 469574 68854 469658
rect 68234 469338 68266 469574
rect 68502 469338 68586 469574
rect 68822 469338 68854 469574
rect 68234 429894 68854 469338
rect 68234 429658 68266 429894
rect 68502 429658 68586 429894
rect 68822 429658 68854 429894
rect 68234 429574 68854 429658
rect 68234 429338 68266 429574
rect 68502 429338 68586 429574
rect 68822 429338 68854 429574
rect 68234 389894 68854 429338
rect 68234 389658 68266 389894
rect 68502 389658 68586 389894
rect 68822 389658 68854 389894
rect 68234 389574 68854 389658
rect 68234 389338 68266 389574
rect 68502 389338 68586 389574
rect 68822 389338 68854 389574
rect 68234 349894 68854 389338
rect 68234 349658 68266 349894
rect 68502 349658 68586 349894
rect 68822 349658 68854 349894
rect 68234 349574 68854 349658
rect 68234 349338 68266 349574
rect 68502 349338 68586 349574
rect 68822 349338 68854 349574
rect 68234 309894 68854 349338
rect 68234 309658 68266 309894
rect 68502 309658 68586 309894
rect 68822 309658 68854 309894
rect 68234 309574 68854 309658
rect 68234 309338 68266 309574
rect 68502 309338 68586 309574
rect 68822 309338 68854 309574
rect 68234 269894 68854 309338
rect 68234 269658 68266 269894
rect 68502 269658 68586 269894
rect 68822 269658 68854 269894
rect 68234 269574 68854 269658
rect 68234 269338 68266 269574
rect 68502 269338 68586 269574
rect 68822 269338 68854 269574
rect 68234 229894 68854 269338
rect 68234 229658 68266 229894
rect 68502 229658 68586 229894
rect 68822 229658 68854 229894
rect 68234 229574 68854 229658
rect 68234 229338 68266 229574
rect 68502 229338 68586 229574
rect 68822 229338 68854 229574
rect 68234 189894 68854 229338
rect 68234 189658 68266 189894
rect 68502 189658 68586 189894
rect 68822 189658 68854 189894
rect 68234 189574 68854 189658
rect 68234 189338 68266 189574
rect 68502 189338 68586 189574
rect 68822 189338 68854 189574
rect 68234 149894 68854 189338
rect 68234 149658 68266 149894
rect 68502 149658 68586 149894
rect 68822 149658 68854 149894
rect 68234 149574 68854 149658
rect 68234 149338 68266 149574
rect 68502 149338 68586 149574
rect 68822 149338 68854 149574
rect 68234 109894 68854 149338
rect 68234 109658 68266 109894
rect 68502 109658 68586 109894
rect 68822 109658 68854 109894
rect 68234 109574 68854 109658
rect 68234 109338 68266 109574
rect 68502 109338 68586 109574
rect 68822 109338 68854 109574
rect 68234 69894 68854 109338
rect 68234 69658 68266 69894
rect 68502 69658 68586 69894
rect 68822 69658 68854 69894
rect 68234 69574 68854 69658
rect 68234 69338 68266 69574
rect 68502 69338 68586 69574
rect 68822 69338 68854 69574
rect 68234 29894 68854 69338
rect 68234 29658 68266 29894
rect 68502 29658 68586 29894
rect 68822 29658 68854 29894
rect 68234 29574 68854 29658
rect 68234 29338 68266 29574
rect 68502 29338 68586 29574
rect 68822 29338 68854 29574
rect 68234 -5146 68854 29338
rect 68234 -5382 68266 -5146
rect 68502 -5382 68586 -5146
rect 68822 -5382 68854 -5146
rect 68234 -5466 68854 -5382
rect 68234 -5702 68266 -5466
rect 68502 -5702 68586 -5466
rect 68822 -5702 68854 -5466
rect 68234 -5734 68854 -5702
rect 71954 673614 72574 711002
rect 91954 710598 92574 711590
rect 91954 710362 91986 710598
rect 92222 710362 92306 710598
rect 92542 710362 92574 710598
rect 91954 710278 92574 710362
rect 91954 710042 91986 710278
rect 92222 710042 92306 710278
rect 92542 710042 92574 710278
rect 88234 708678 88854 709670
rect 88234 708442 88266 708678
rect 88502 708442 88586 708678
rect 88822 708442 88854 708678
rect 88234 708358 88854 708442
rect 88234 708122 88266 708358
rect 88502 708122 88586 708358
rect 88822 708122 88854 708358
rect 84514 706758 85134 707750
rect 84514 706522 84546 706758
rect 84782 706522 84866 706758
rect 85102 706522 85134 706758
rect 84514 706438 85134 706522
rect 84514 706202 84546 706438
rect 84782 706202 84866 706438
rect 85102 706202 85134 706438
rect 71954 673378 71986 673614
rect 72222 673378 72306 673614
rect 72542 673378 72574 673614
rect 71954 673294 72574 673378
rect 71954 673058 71986 673294
rect 72222 673058 72306 673294
rect 72542 673058 72574 673294
rect 71954 633614 72574 673058
rect 71954 633378 71986 633614
rect 72222 633378 72306 633614
rect 72542 633378 72574 633614
rect 71954 633294 72574 633378
rect 71954 633058 71986 633294
rect 72222 633058 72306 633294
rect 72542 633058 72574 633294
rect 71954 593614 72574 633058
rect 71954 593378 71986 593614
rect 72222 593378 72306 593614
rect 72542 593378 72574 593614
rect 71954 593294 72574 593378
rect 71954 593058 71986 593294
rect 72222 593058 72306 593294
rect 72542 593058 72574 593294
rect 71954 553614 72574 593058
rect 71954 553378 71986 553614
rect 72222 553378 72306 553614
rect 72542 553378 72574 553614
rect 71954 553294 72574 553378
rect 71954 553058 71986 553294
rect 72222 553058 72306 553294
rect 72542 553058 72574 553294
rect 71954 513614 72574 553058
rect 71954 513378 71986 513614
rect 72222 513378 72306 513614
rect 72542 513378 72574 513614
rect 71954 513294 72574 513378
rect 71954 513058 71986 513294
rect 72222 513058 72306 513294
rect 72542 513058 72574 513294
rect 71954 473614 72574 513058
rect 71954 473378 71986 473614
rect 72222 473378 72306 473614
rect 72542 473378 72574 473614
rect 71954 473294 72574 473378
rect 71954 473058 71986 473294
rect 72222 473058 72306 473294
rect 72542 473058 72574 473294
rect 71954 433614 72574 473058
rect 71954 433378 71986 433614
rect 72222 433378 72306 433614
rect 72542 433378 72574 433614
rect 71954 433294 72574 433378
rect 71954 433058 71986 433294
rect 72222 433058 72306 433294
rect 72542 433058 72574 433294
rect 71954 393614 72574 433058
rect 71954 393378 71986 393614
rect 72222 393378 72306 393614
rect 72542 393378 72574 393614
rect 71954 393294 72574 393378
rect 71954 393058 71986 393294
rect 72222 393058 72306 393294
rect 72542 393058 72574 393294
rect 71954 353614 72574 393058
rect 71954 353378 71986 353614
rect 72222 353378 72306 353614
rect 72542 353378 72574 353614
rect 71954 353294 72574 353378
rect 71954 353058 71986 353294
rect 72222 353058 72306 353294
rect 72542 353058 72574 353294
rect 71954 313614 72574 353058
rect 71954 313378 71986 313614
rect 72222 313378 72306 313614
rect 72542 313378 72574 313614
rect 71954 313294 72574 313378
rect 71954 313058 71986 313294
rect 72222 313058 72306 313294
rect 72542 313058 72574 313294
rect 71954 273614 72574 313058
rect 71954 273378 71986 273614
rect 72222 273378 72306 273614
rect 72542 273378 72574 273614
rect 71954 273294 72574 273378
rect 71954 273058 71986 273294
rect 72222 273058 72306 273294
rect 72542 273058 72574 273294
rect 71954 233614 72574 273058
rect 71954 233378 71986 233614
rect 72222 233378 72306 233614
rect 72542 233378 72574 233614
rect 71954 233294 72574 233378
rect 71954 233058 71986 233294
rect 72222 233058 72306 233294
rect 72542 233058 72574 233294
rect 71954 193614 72574 233058
rect 71954 193378 71986 193614
rect 72222 193378 72306 193614
rect 72542 193378 72574 193614
rect 71954 193294 72574 193378
rect 71954 193058 71986 193294
rect 72222 193058 72306 193294
rect 72542 193058 72574 193294
rect 71954 153614 72574 193058
rect 71954 153378 71986 153614
rect 72222 153378 72306 153614
rect 72542 153378 72574 153614
rect 71954 153294 72574 153378
rect 71954 153058 71986 153294
rect 72222 153058 72306 153294
rect 72542 153058 72574 153294
rect 71954 113614 72574 153058
rect 71954 113378 71986 113614
rect 72222 113378 72306 113614
rect 72542 113378 72574 113614
rect 71954 113294 72574 113378
rect 71954 113058 71986 113294
rect 72222 113058 72306 113294
rect 72542 113058 72574 113294
rect 71954 73614 72574 113058
rect 71954 73378 71986 73614
rect 72222 73378 72306 73614
rect 72542 73378 72574 73614
rect 71954 73294 72574 73378
rect 71954 73058 71986 73294
rect 72222 73058 72306 73294
rect 72542 73058 72574 73294
rect 71954 33614 72574 73058
rect 71954 33378 71986 33614
rect 72222 33378 72306 33614
rect 72542 33378 72574 33614
rect 71954 33294 72574 33378
rect 71954 33058 71986 33294
rect 72222 33058 72306 33294
rect 72542 33058 72574 33294
rect 51954 -6342 51986 -6106
rect 52222 -6342 52306 -6106
rect 52542 -6342 52574 -6106
rect 51954 -6426 52574 -6342
rect 51954 -6662 51986 -6426
rect 52222 -6662 52306 -6426
rect 52542 -6662 52574 -6426
rect 51954 -7654 52574 -6662
rect 71954 -7066 72574 33058
rect 80794 704838 81414 705830
rect 80794 704602 80826 704838
rect 81062 704602 81146 704838
rect 81382 704602 81414 704838
rect 80794 704518 81414 704602
rect 80794 704282 80826 704518
rect 81062 704282 81146 704518
rect 81382 704282 81414 704518
rect 80794 682454 81414 704282
rect 80794 682218 80826 682454
rect 81062 682218 81146 682454
rect 81382 682218 81414 682454
rect 80794 682134 81414 682218
rect 80794 681898 80826 682134
rect 81062 681898 81146 682134
rect 81382 681898 81414 682134
rect 80794 642454 81414 681898
rect 80794 642218 80826 642454
rect 81062 642218 81146 642454
rect 81382 642218 81414 642454
rect 80794 642134 81414 642218
rect 80794 641898 80826 642134
rect 81062 641898 81146 642134
rect 81382 641898 81414 642134
rect 80794 602454 81414 641898
rect 80794 602218 80826 602454
rect 81062 602218 81146 602454
rect 81382 602218 81414 602454
rect 80794 602134 81414 602218
rect 80794 601898 80826 602134
rect 81062 601898 81146 602134
rect 81382 601898 81414 602134
rect 80794 562454 81414 601898
rect 80794 562218 80826 562454
rect 81062 562218 81146 562454
rect 81382 562218 81414 562454
rect 80794 562134 81414 562218
rect 80794 561898 80826 562134
rect 81062 561898 81146 562134
rect 81382 561898 81414 562134
rect 80794 522454 81414 561898
rect 80794 522218 80826 522454
rect 81062 522218 81146 522454
rect 81382 522218 81414 522454
rect 80794 522134 81414 522218
rect 80794 521898 80826 522134
rect 81062 521898 81146 522134
rect 81382 521898 81414 522134
rect 80794 482454 81414 521898
rect 80794 482218 80826 482454
rect 81062 482218 81146 482454
rect 81382 482218 81414 482454
rect 80794 482134 81414 482218
rect 80794 481898 80826 482134
rect 81062 481898 81146 482134
rect 81382 481898 81414 482134
rect 80794 442454 81414 481898
rect 80794 442218 80826 442454
rect 81062 442218 81146 442454
rect 81382 442218 81414 442454
rect 80794 442134 81414 442218
rect 80794 441898 80826 442134
rect 81062 441898 81146 442134
rect 81382 441898 81414 442134
rect 80794 402454 81414 441898
rect 80794 402218 80826 402454
rect 81062 402218 81146 402454
rect 81382 402218 81414 402454
rect 80794 402134 81414 402218
rect 80794 401898 80826 402134
rect 81062 401898 81146 402134
rect 81382 401898 81414 402134
rect 80794 362454 81414 401898
rect 80794 362218 80826 362454
rect 81062 362218 81146 362454
rect 81382 362218 81414 362454
rect 80794 362134 81414 362218
rect 80794 361898 80826 362134
rect 81062 361898 81146 362134
rect 81382 361898 81414 362134
rect 80794 322454 81414 361898
rect 80794 322218 80826 322454
rect 81062 322218 81146 322454
rect 81382 322218 81414 322454
rect 80794 322134 81414 322218
rect 80794 321898 80826 322134
rect 81062 321898 81146 322134
rect 81382 321898 81414 322134
rect 80794 282454 81414 321898
rect 80794 282218 80826 282454
rect 81062 282218 81146 282454
rect 81382 282218 81414 282454
rect 80794 282134 81414 282218
rect 80794 281898 80826 282134
rect 81062 281898 81146 282134
rect 81382 281898 81414 282134
rect 80794 242454 81414 281898
rect 80794 242218 80826 242454
rect 81062 242218 81146 242454
rect 81382 242218 81414 242454
rect 80794 242134 81414 242218
rect 80794 241898 80826 242134
rect 81062 241898 81146 242134
rect 81382 241898 81414 242134
rect 80794 202454 81414 241898
rect 80794 202218 80826 202454
rect 81062 202218 81146 202454
rect 81382 202218 81414 202454
rect 80794 202134 81414 202218
rect 80794 201898 80826 202134
rect 81062 201898 81146 202134
rect 81382 201898 81414 202134
rect 80794 162454 81414 201898
rect 80794 162218 80826 162454
rect 81062 162218 81146 162454
rect 81382 162218 81414 162454
rect 80794 162134 81414 162218
rect 80794 161898 80826 162134
rect 81062 161898 81146 162134
rect 81382 161898 81414 162134
rect 80794 122454 81414 161898
rect 80794 122218 80826 122454
rect 81062 122218 81146 122454
rect 81382 122218 81414 122454
rect 80794 122134 81414 122218
rect 80794 121898 80826 122134
rect 81062 121898 81146 122134
rect 81382 121898 81414 122134
rect 80794 82454 81414 121898
rect 80794 82218 80826 82454
rect 81062 82218 81146 82454
rect 81382 82218 81414 82454
rect 80794 82134 81414 82218
rect 80794 81898 80826 82134
rect 81062 81898 81146 82134
rect 81382 81898 81414 82134
rect 80794 42454 81414 81898
rect 80794 42218 80826 42454
rect 81062 42218 81146 42454
rect 81382 42218 81414 42454
rect 80794 42134 81414 42218
rect 80794 41898 80826 42134
rect 81062 41898 81146 42134
rect 81382 41898 81414 42134
rect 80794 2454 81414 41898
rect 80794 2218 80826 2454
rect 81062 2218 81146 2454
rect 81382 2218 81414 2454
rect 80794 2134 81414 2218
rect 80794 1898 80826 2134
rect 81062 1898 81146 2134
rect 81382 1898 81414 2134
rect 80794 -346 81414 1898
rect 80794 -582 80826 -346
rect 81062 -582 81146 -346
rect 81382 -582 81414 -346
rect 80794 -666 81414 -582
rect 80794 -902 80826 -666
rect 81062 -902 81146 -666
rect 81382 -902 81414 -666
rect 80794 -1894 81414 -902
rect 84514 686174 85134 706202
rect 84514 685938 84546 686174
rect 84782 685938 84866 686174
rect 85102 685938 85134 686174
rect 84514 685854 85134 685938
rect 84514 685618 84546 685854
rect 84782 685618 84866 685854
rect 85102 685618 85134 685854
rect 84514 646174 85134 685618
rect 84514 645938 84546 646174
rect 84782 645938 84866 646174
rect 85102 645938 85134 646174
rect 84514 645854 85134 645938
rect 84514 645618 84546 645854
rect 84782 645618 84866 645854
rect 85102 645618 85134 645854
rect 84514 606174 85134 645618
rect 84514 605938 84546 606174
rect 84782 605938 84866 606174
rect 85102 605938 85134 606174
rect 84514 605854 85134 605938
rect 84514 605618 84546 605854
rect 84782 605618 84866 605854
rect 85102 605618 85134 605854
rect 84514 566174 85134 605618
rect 84514 565938 84546 566174
rect 84782 565938 84866 566174
rect 85102 565938 85134 566174
rect 84514 565854 85134 565938
rect 84514 565618 84546 565854
rect 84782 565618 84866 565854
rect 85102 565618 85134 565854
rect 84514 526174 85134 565618
rect 84514 525938 84546 526174
rect 84782 525938 84866 526174
rect 85102 525938 85134 526174
rect 84514 525854 85134 525938
rect 84514 525618 84546 525854
rect 84782 525618 84866 525854
rect 85102 525618 85134 525854
rect 84514 486174 85134 525618
rect 84514 485938 84546 486174
rect 84782 485938 84866 486174
rect 85102 485938 85134 486174
rect 84514 485854 85134 485938
rect 84514 485618 84546 485854
rect 84782 485618 84866 485854
rect 85102 485618 85134 485854
rect 84514 446174 85134 485618
rect 84514 445938 84546 446174
rect 84782 445938 84866 446174
rect 85102 445938 85134 446174
rect 84514 445854 85134 445938
rect 84514 445618 84546 445854
rect 84782 445618 84866 445854
rect 85102 445618 85134 445854
rect 84514 406174 85134 445618
rect 84514 405938 84546 406174
rect 84782 405938 84866 406174
rect 85102 405938 85134 406174
rect 84514 405854 85134 405938
rect 84514 405618 84546 405854
rect 84782 405618 84866 405854
rect 85102 405618 85134 405854
rect 84514 366174 85134 405618
rect 84514 365938 84546 366174
rect 84782 365938 84866 366174
rect 85102 365938 85134 366174
rect 84514 365854 85134 365938
rect 84514 365618 84546 365854
rect 84782 365618 84866 365854
rect 85102 365618 85134 365854
rect 84514 326174 85134 365618
rect 84514 325938 84546 326174
rect 84782 325938 84866 326174
rect 85102 325938 85134 326174
rect 84514 325854 85134 325938
rect 84514 325618 84546 325854
rect 84782 325618 84866 325854
rect 85102 325618 85134 325854
rect 84514 286174 85134 325618
rect 84514 285938 84546 286174
rect 84782 285938 84866 286174
rect 85102 285938 85134 286174
rect 84514 285854 85134 285938
rect 84514 285618 84546 285854
rect 84782 285618 84866 285854
rect 85102 285618 85134 285854
rect 84514 246174 85134 285618
rect 84514 245938 84546 246174
rect 84782 245938 84866 246174
rect 85102 245938 85134 246174
rect 84514 245854 85134 245938
rect 84514 245618 84546 245854
rect 84782 245618 84866 245854
rect 85102 245618 85134 245854
rect 84514 206174 85134 245618
rect 84514 205938 84546 206174
rect 84782 205938 84866 206174
rect 85102 205938 85134 206174
rect 84514 205854 85134 205938
rect 84514 205618 84546 205854
rect 84782 205618 84866 205854
rect 85102 205618 85134 205854
rect 84514 166174 85134 205618
rect 84514 165938 84546 166174
rect 84782 165938 84866 166174
rect 85102 165938 85134 166174
rect 84514 165854 85134 165938
rect 84514 165618 84546 165854
rect 84782 165618 84866 165854
rect 85102 165618 85134 165854
rect 84514 126174 85134 165618
rect 84514 125938 84546 126174
rect 84782 125938 84866 126174
rect 85102 125938 85134 126174
rect 84514 125854 85134 125938
rect 84514 125618 84546 125854
rect 84782 125618 84866 125854
rect 85102 125618 85134 125854
rect 84514 86174 85134 125618
rect 84514 85938 84546 86174
rect 84782 85938 84866 86174
rect 85102 85938 85134 86174
rect 84514 85854 85134 85938
rect 84514 85618 84546 85854
rect 84782 85618 84866 85854
rect 85102 85618 85134 85854
rect 84514 46174 85134 85618
rect 84514 45938 84546 46174
rect 84782 45938 84866 46174
rect 85102 45938 85134 46174
rect 84514 45854 85134 45938
rect 84514 45618 84546 45854
rect 84782 45618 84866 45854
rect 85102 45618 85134 45854
rect 84514 6174 85134 45618
rect 84514 5938 84546 6174
rect 84782 5938 84866 6174
rect 85102 5938 85134 6174
rect 84514 5854 85134 5938
rect 84514 5618 84546 5854
rect 84782 5618 84866 5854
rect 85102 5618 85134 5854
rect 84514 -2266 85134 5618
rect 84514 -2502 84546 -2266
rect 84782 -2502 84866 -2266
rect 85102 -2502 85134 -2266
rect 84514 -2586 85134 -2502
rect 84514 -2822 84546 -2586
rect 84782 -2822 84866 -2586
rect 85102 -2822 85134 -2586
rect 84514 -3814 85134 -2822
rect 88234 689894 88854 708122
rect 88234 689658 88266 689894
rect 88502 689658 88586 689894
rect 88822 689658 88854 689894
rect 88234 689574 88854 689658
rect 88234 689338 88266 689574
rect 88502 689338 88586 689574
rect 88822 689338 88854 689574
rect 88234 649894 88854 689338
rect 88234 649658 88266 649894
rect 88502 649658 88586 649894
rect 88822 649658 88854 649894
rect 88234 649574 88854 649658
rect 88234 649338 88266 649574
rect 88502 649338 88586 649574
rect 88822 649338 88854 649574
rect 88234 609894 88854 649338
rect 88234 609658 88266 609894
rect 88502 609658 88586 609894
rect 88822 609658 88854 609894
rect 88234 609574 88854 609658
rect 88234 609338 88266 609574
rect 88502 609338 88586 609574
rect 88822 609338 88854 609574
rect 88234 569894 88854 609338
rect 88234 569658 88266 569894
rect 88502 569658 88586 569894
rect 88822 569658 88854 569894
rect 88234 569574 88854 569658
rect 88234 569338 88266 569574
rect 88502 569338 88586 569574
rect 88822 569338 88854 569574
rect 88234 529894 88854 569338
rect 88234 529658 88266 529894
rect 88502 529658 88586 529894
rect 88822 529658 88854 529894
rect 88234 529574 88854 529658
rect 88234 529338 88266 529574
rect 88502 529338 88586 529574
rect 88822 529338 88854 529574
rect 88234 489894 88854 529338
rect 88234 489658 88266 489894
rect 88502 489658 88586 489894
rect 88822 489658 88854 489894
rect 88234 489574 88854 489658
rect 88234 489338 88266 489574
rect 88502 489338 88586 489574
rect 88822 489338 88854 489574
rect 88234 449894 88854 489338
rect 88234 449658 88266 449894
rect 88502 449658 88586 449894
rect 88822 449658 88854 449894
rect 88234 449574 88854 449658
rect 88234 449338 88266 449574
rect 88502 449338 88586 449574
rect 88822 449338 88854 449574
rect 88234 409894 88854 449338
rect 88234 409658 88266 409894
rect 88502 409658 88586 409894
rect 88822 409658 88854 409894
rect 88234 409574 88854 409658
rect 88234 409338 88266 409574
rect 88502 409338 88586 409574
rect 88822 409338 88854 409574
rect 88234 369894 88854 409338
rect 88234 369658 88266 369894
rect 88502 369658 88586 369894
rect 88822 369658 88854 369894
rect 88234 369574 88854 369658
rect 88234 369338 88266 369574
rect 88502 369338 88586 369574
rect 88822 369338 88854 369574
rect 88234 329894 88854 369338
rect 88234 329658 88266 329894
rect 88502 329658 88586 329894
rect 88822 329658 88854 329894
rect 88234 329574 88854 329658
rect 88234 329338 88266 329574
rect 88502 329338 88586 329574
rect 88822 329338 88854 329574
rect 88234 289894 88854 329338
rect 88234 289658 88266 289894
rect 88502 289658 88586 289894
rect 88822 289658 88854 289894
rect 88234 289574 88854 289658
rect 88234 289338 88266 289574
rect 88502 289338 88586 289574
rect 88822 289338 88854 289574
rect 88234 249894 88854 289338
rect 88234 249658 88266 249894
rect 88502 249658 88586 249894
rect 88822 249658 88854 249894
rect 88234 249574 88854 249658
rect 88234 249338 88266 249574
rect 88502 249338 88586 249574
rect 88822 249338 88854 249574
rect 88234 209894 88854 249338
rect 88234 209658 88266 209894
rect 88502 209658 88586 209894
rect 88822 209658 88854 209894
rect 88234 209574 88854 209658
rect 88234 209338 88266 209574
rect 88502 209338 88586 209574
rect 88822 209338 88854 209574
rect 88234 169894 88854 209338
rect 88234 169658 88266 169894
rect 88502 169658 88586 169894
rect 88822 169658 88854 169894
rect 88234 169574 88854 169658
rect 88234 169338 88266 169574
rect 88502 169338 88586 169574
rect 88822 169338 88854 169574
rect 88234 129894 88854 169338
rect 88234 129658 88266 129894
rect 88502 129658 88586 129894
rect 88822 129658 88854 129894
rect 88234 129574 88854 129658
rect 88234 129338 88266 129574
rect 88502 129338 88586 129574
rect 88822 129338 88854 129574
rect 88234 89894 88854 129338
rect 88234 89658 88266 89894
rect 88502 89658 88586 89894
rect 88822 89658 88854 89894
rect 88234 89574 88854 89658
rect 88234 89338 88266 89574
rect 88502 89338 88586 89574
rect 88822 89338 88854 89574
rect 88234 49894 88854 89338
rect 88234 49658 88266 49894
rect 88502 49658 88586 49894
rect 88822 49658 88854 49894
rect 88234 49574 88854 49658
rect 88234 49338 88266 49574
rect 88502 49338 88586 49574
rect 88822 49338 88854 49574
rect 88234 9894 88854 49338
rect 88234 9658 88266 9894
rect 88502 9658 88586 9894
rect 88822 9658 88854 9894
rect 88234 9574 88854 9658
rect 88234 9338 88266 9574
rect 88502 9338 88586 9574
rect 88822 9338 88854 9574
rect 88234 -4186 88854 9338
rect 88234 -4422 88266 -4186
rect 88502 -4422 88586 -4186
rect 88822 -4422 88854 -4186
rect 88234 -4506 88854 -4422
rect 88234 -4742 88266 -4506
rect 88502 -4742 88586 -4506
rect 88822 -4742 88854 -4506
rect 88234 -5734 88854 -4742
rect 91954 693614 92574 710042
rect 111954 711558 112574 711590
rect 111954 711322 111986 711558
rect 112222 711322 112306 711558
rect 112542 711322 112574 711558
rect 111954 711238 112574 711322
rect 111954 711002 111986 711238
rect 112222 711002 112306 711238
rect 112542 711002 112574 711238
rect 108234 709638 108854 709670
rect 108234 709402 108266 709638
rect 108502 709402 108586 709638
rect 108822 709402 108854 709638
rect 108234 709318 108854 709402
rect 108234 709082 108266 709318
rect 108502 709082 108586 709318
rect 108822 709082 108854 709318
rect 104514 707718 105134 707750
rect 104514 707482 104546 707718
rect 104782 707482 104866 707718
rect 105102 707482 105134 707718
rect 104514 707398 105134 707482
rect 104514 707162 104546 707398
rect 104782 707162 104866 707398
rect 105102 707162 105134 707398
rect 91954 693378 91986 693614
rect 92222 693378 92306 693614
rect 92542 693378 92574 693614
rect 91954 693294 92574 693378
rect 91954 693058 91986 693294
rect 92222 693058 92306 693294
rect 92542 693058 92574 693294
rect 91954 653614 92574 693058
rect 91954 653378 91986 653614
rect 92222 653378 92306 653614
rect 92542 653378 92574 653614
rect 91954 653294 92574 653378
rect 91954 653058 91986 653294
rect 92222 653058 92306 653294
rect 92542 653058 92574 653294
rect 91954 613614 92574 653058
rect 91954 613378 91986 613614
rect 92222 613378 92306 613614
rect 92542 613378 92574 613614
rect 91954 613294 92574 613378
rect 91954 613058 91986 613294
rect 92222 613058 92306 613294
rect 92542 613058 92574 613294
rect 91954 573614 92574 613058
rect 91954 573378 91986 573614
rect 92222 573378 92306 573614
rect 92542 573378 92574 573614
rect 91954 573294 92574 573378
rect 91954 573058 91986 573294
rect 92222 573058 92306 573294
rect 92542 573058 92574 573294
rect 91954 533614 92574 573058
rect 91954 533378 91986 533614
rect 92222 533378 92306 533614
rect 92542 533378 92574 533614
rect 91954 533294 92574 533378
rect 91954 533058 91986 533294
rect 92222 533058 92306 533294
rect 92542 533058 92574 533294
rect 91954 493614 92574 533058
rect 91954 493378 91986 493614
rect 92222 493378 92306 493614
rect 92542 493378 92574 493614
rect 91954 493294 92574 493378
rect 91954 493058 91986 493294
rect 92222 493058 92306 493294
rect 92542 493058 92574 493294
rect 91954 453614 92574 493058
rect 91954 453378 91986 453614
rect 92222 453378 92306 453614
rect 92542 453378 92574 453614
rect 91954 453294 92574 453378
rect 91954 453058 91986 453294
rect 92222 453058 92306 453294
rect 92542 453058 92574 453294
rect 91954 413614 92574 453058
rect 91954 413378 91986 413614
rect 92222 413378 92306 413614
rect 92542 413378 92574 413614
rect 91954 413294 92574 413378
rect 91954 413058 91986 413294
rect 92222 413058 92306 413294
rect 92542 413058 92574 413294
rect 91954 373614 92574 413058
rect 91954 373378 91986 373614
rect 92222 373378 92306 373614
rect 92542 373378 92574 373614
rect 91954 373294 92574 373378
rect 91954 373058 91986 373294
rect 92222 373058 92306 373294
rect 92542 373058 92574 373294
rect 91954 333614 92574 373058
rect 91954 333378 91986 333614
rect 92222 333378 92306 333614
rect 92542 333378 92574 333614
rect 91954 333294 92574 333378
rect 91954 333058 91986 333294
rect 92222 333058 92306 333294
rect 92542 333058 92574 333294
rect 91954 293614 92574 333058
rect 91954 293378 91986 293614
rect 92222 293378 92306 293614
rect 92542 293378 92574 293614
rect 91954 293294 92574 293378
rect 91954 293058 91986 293294
rect 92222 293058 92306 293294
rect 92542 293058 92574 293294
rect 91954 253614 92574 293058
rect 91954 253378 91986 253614
rect 92222 253378 92306 253614
rect 92542 253378 92574 253614
rect 91954 253294 92574 253378
rect 91954 253058 91986 253294
rect 92222 253058 92306 253294
rect 92542 253058 92574 253294
rect 91954 213614 92574 253058
rect 91954 213378 91986 213614
rect 92222 213378 92306 213614
rect 92542 213378 92574 213614
rect 91954 213294 92574 213378
rect 91954 213058 91986 213294
rect 92222 213058 92306 213294
rect 92542 213058 92574 213294
rect 91954 173614 92574 213058
rect 91954 173378 91986 173614
rect 92222 173378 92306 173614
rect 92542 173378 92574 173614
rect 91954 173294 92574 173378
rect 91954 173058 91986 173294
rect 92222 173058 92306 173294
rect 92542 173058 92574 173294
rect 91954 133614 92574 173058
rect 91954 133378 91986 133614
rect 92222 133378 92306 133614
rect 92542 133378 92574 133614
rect 91954 133294 92574 133378
rect 91954 133058 91986 133294
rect 92222 133058 92306 133294
rect 92542 133058 92574 133294
rect 91954 93614 92574 133058
rect 91954 93378 91986 93614
rect 92222 93378 92306 93614
rect 92542 93378 92574 93614
rect 91954 93294 92574 93378
rect 91954 93058 91986 93294
rect 92222 93058 92306 93294
rect 92542 93058 92574 93294
rect 91954 53614 92574 93058
rect 91954 53378 91986 53614
rect 92222 53378 92306 53614
rect 92542 53378 92574 53614
rect 91954 53294 92574 53378
rect 91954 53058 91986 53294
rect 92222 53058 92306 53294
rect 92542 53058 92574 53294
rect 91954 13614 92574 53058
rect 91954 13378 91986 13614
rect 92222 13378 92306 13614
rect 92542 13378 92574 13614
rect 91954 13294 92574 13378
rect 91954 13058 91986 13294
rect 92222 13058 92306 13294
rect 92542 13058 92574 13294
rect 71954 -7302 71986 -7066
rect 72222 -7302 72306 -7066
rect 72542 -7302 72574 -7066
rect 71954 -7386 72574 -7302
rect 71954 -7622 71986 -7386
rect 72222 -7622 72306 -7386
rect 72542 -7622 72574 -7386
rect 71954 -7654 72574 -7622
rect 91954 -6106 92574 13058
rect 100794 705798 101414 705830
rect 100794 705562 100826 705798
rect 101062 705562 101146 705798
rect 101382 705562 101414 705798
rect 100794 705478 101414 705562
rect 100794 705242 100826 705478
rect 101062 705242 101146 705478
rect 101382 705242 101414 705478
rect 100794 662454 101414 705242
rect 100794 662218 100826 662454
rect 101062 662218 101146 662454
rect 101382 662218 101414 662454
rect 100794 662134 101414 662218
rect 100794 661898 100826 662134
rect 101062 661898 101146 662134
rect 101382 661898 101414 662134
rect 100794 622454 101414 661898
rect 100794 622218 100826 622454
rect 101062 622218 101146 622454
rect 101382 622218 101414 622454
rect 100794 622134 101414 622218
rect 100794 621898 100826 622134
rect 101062 621898 101146 622134
rect 101382 621898 101414 622134
rect 100794 582454 101414 621898
rect 100794 582218 100826 582454
rect 101062 582218 101146 582454
rect 101382 582218 101414 582454
rect 100794 582134 101414 582218
rect 100794 581898 100826 582134
rect 101062 581898 101146 582134
rect 101382 581898 101414 582134
rect 100794 542454 101414 581898
rect 100794 542218 100826 542454
rect 101062 542218 101146 542454
rect 101382 542218 101414 542454
rect 100794 542134 101414 542218
rect 100794 541898 100826 542134
rect 101062 541898 101146 542134
rect 101382 541898 101414 542134
rect 100794 502454 101414 541898
rect 100794 502218 100826 502454
rect 101062 502218 101146 502454
rect 101382 502218 101414 502454
rect 100794 502134 101414 502218
rect 100794 501898 100826 502134
rect 101062 501898 101146 502134
rect 101382 501898 101414 502134
rect 100794 462454 101414 501898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 422454 101414 461898
rect 100794 422218 100826 422454
rect 101062 422218 101146 422454
rect 101382 422218 101414 422454
rect 100794 422134 101414 422218
rect 100794 421898 100826 422134
rect 101062 421898 101146 422134
rect 101382 421898 101414 422134
rect 100794 382454 101414 421898
rect 100794 382218 100826 382454
rect 101062 382218 101146 382454
rect 101382 382218 101414 382454
rect 100794 382134 101414 382218
rect 100794 381898 100826 382134
rect 101062 381898 101146 382134
rect 101382 381898 101414 382134
rect 100794 342454 101414 381898
rect 100794 342218 100826 342454
rect 101062 342218 101146 342454
rect 101382 342218 101414 342454
rect 100794 342134 101414 342218
rect 100794 341898 100826 342134
rect 101062 341898 101146 342134
rect 101382 341898 101414 342134
rect 100794 302454 101414 341898
rect 100794 302218 100826 302454
rect 101062 302218 101146 302454
rect 101382 302218 101414 302454
rect 100794 302134 101414 302218
rect 100794 301898 100826 302134
rect 101062 301898 101146 302134
rect 101382 301898 101414 302134
rect 100794 262454 101414 301898
rect 100794 262218 100826 262454
rect 101062 262218 101146 262454
rect 101382 262218 101414 262454
rect 100794 262134 101414 262218
rect 100794 261898 100826 262134
rect 101062 261898 101146 262134
rect 101382 261898 101414 262134
rect 100794 222454 101414 261898
rect 100794 222218 100826 222454
rect 101062 222218 101146 222454
rect 101382 222218 101414 222454
rect 100794 222134 101414 222218
rect 100794 221898 100826 222134
rect 101062 221898 101146 222134
rect 101382 221898 101414 222134
rect 100794 182454 101414 221898
rect 100794 182218 100826 182454
rect 101062 182218 101146 182454
rect 101382 182218 101414 182454
rect 100794 182134 101414 182218
rect 100794 181898 100826 182134
rect 101062 181898 101146 182134
rect 101382 181898 101414 182134
rect 100794 142454 101414 181898
rect 100794 142218 100826 142454
rect 101062 142218 101146 142454
rect 101382 142218 101414 142454
rect 100794 142134 101414 142218
rect 100794 141898 100826 142134
rect 101062 141898 101146 142134
rect 101382 141898 101414 142134
rect 100794 102454 101414 141898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 62454 101414 101898
rect 100794 62218 100826 62454
rect 101062 62218 101146 62454
rect 101382 62218 101414 62454
rect 100794 62134 101414 62218
rect 100794 61898 100826 62134
rect 101062 61898 101146 62134
rect 101382 61898 101414 62134
rect 100794 22454 101414 61898
rect 100794 22218 100826 22454
rect 101062 22218 101146 22454
rect 101382 22218 101414 22454
rect 100794 22134 101414 22218
rect 100794 21898 100826 22134
rect 101062 21898 101146 22134
rect 101382 21898 101414 22134
rect 100794 -1306 101414 21898
rect 100794 -1542 100826 -1306
rect 101062 -1542 101146 -1306
rect 101382 -1542 101414 -1306
rect 100794 -1626 101414 -1542
rect 100794 -1862 100826 -1626
rect 101062 -1862 101146 -1626
rect 101382 -1862 101414 -1626
rect 100794 -1894 101414 -1862
rect 104514 666174 105134 707162
rect 104514 665938 104546 666174
rect 104782 665938 104866 666174
rect 105102 665938 105134 666174
rect 104514 665854 105134 665938
rect 104514 665618 104546 665854
rect 104782 665618 104866 665854
rect 105102 665618 105134 665854
rect 104514 626174 105134 665618
rect 104514 625938 104546 626174
rect 104782 625938 104866 626174
rect 105102 625938 105134 626174
rect 104514 625854 105134 625938
rect 104514 625618 104546 625854
rect 104782 625618 104866 625854
rect 105102 625618 105134 625854
rect 104514 586174 105134 625618
rect 104514 585938 104546 586174
rect 104782 585938 104866 586174
rect 105102 585938 105134 586174
rect 104514 585854 105134 585938
rect 104514 585618 104546 585854
rect 104782 585618 104866 585854
rect 105102 585618 105134 585854
rect 104514 546174 105134 585618
rect 104514 545938 104546 546174
rect 104782 545938 104866 546174
rect 105102 545938 105134 546174
rect 104514 545854 105134 545938
rect 104514 545618 104546 545854
rect 104782 545618 104866 545854
rect 105102 545618 105134 545854
rect 104514 506174 105134 545618
rect 104514 505938 104546 506174
rect 104782 505938 104866 506174
rect 105102 505938 105134 506174
rect 104514 505854 105134 505938
rect 104514 505618 104546 505854
rect 104782 505618 104866 505854
rect 105102 505618 105134 505854
rect 104514 466174 105134 505618
rect 104514 465938 104546 466174
rect 104782 465938 104866 466174
rect 105102 465938 105134 466174
rect 104514 465854 105134 465938
rect 104514 465618 104546 465854
rect 104782 465618 104866 465854
rect 105102 465618 105134 465854
rect 104514 426174 105134 465618
rect 104514 425938 104546 426174
rect 104782 425938 104866 426174
rect 105102 425938 105134 426174
rect 104514 425854 105134 425938
rect 104514 425618 104546 425854
rect 104782 425618 104866 425854
rect 105102 425618 105134 425854
rect 104514 386174 105134 425618
rect 104514 385938 104546 386174
rect 104782 385938 104866 386174
rect 105102 385938 105134 386174
rect 104514 385854 105134 385938
rect 104514 385618 104546 385854
rect 104782 385618 104866 385854
rect 105102 385618 105134 385854
rect 104514 346174 105134 385618
rect 104514 345938 104546 346174
rect 104782 345938 104866 346174
rect 105102 345938 105134 346174
rect 104514 345854 105134 345938
rect 104514 345618 104546 345854
rect 104782 345618 104866 345854
rect 105102 345618 105134 345854
rect 104514 306174 105134 345618
rect 104514 305938 104546 306174
rect 104782 305938 104866 306174
rect 105102 305938 105134 306174
rect 104514 305854 105134 305938
rect 104514 305618 104546 305854
rect 104782 305618 104866 305854
rect 105102 305618 105134 305854
rect 104514 266174 105134 305618
rect 104514 265938 104546 266174
rect 104782 265938 104866 266174
rect 105102 265938 105134 266174
rect 104514 265854 105134 265938
rect 104514 265618 104546 265854
rect 104782 265618 104866 265854
rect 105102 265618 105134 265854
rect 104514 226174 105134 265618
rect 104514 225938 104546 226174
rect 104782 225938 104866 226174
rect 105102 225938 105134 226174
rect 104514 225854 105134 225938
rect 104514 225618 104546 225854
rect 104782 225618 104866 225854
rect 105102 225618 105134 225854
rect 104514 186174 105134 225618
rect 104514 185938 104546 186174
rect 104782 185938 104866 186174
rect 105102 185938 105134 186174
rect 104514 185854 105134 185938
rect 104514 185618 104546 185854
rect 104782 185618 104866 185854
rect 105102 185618 105134 185854
rect 104514 146174 105134 185618
rect 104514 145938 104546 146174
rect 104782 145938 104866 146174
rect 105102 145938 105134 146174
rect 104514 145854 105134 145938
rect 104514 145618 104546 145854
rect 104782 145618 104866 145854
rect 105102 145618 105134 145854
rect 104514 106174 105134 145618
rect 104514 105938 104546 106174
rect 104782 105938 104866 106174
rect 105102 105938 105134 106174
rect 104514 105854 105134 105938
rect 104514 105618 104546 105854
rect 104782 105618 104866 105854
rect 105102 105618 105134 105854
rect 104514 66174 105134 105618
rect 104514 65938 104546 66174
rect 104782 65938 104866 66174
rect 105102 65938 105134 66174
rect 104514 65854 105134 65938
rect 104514 65618 104546 65854
rect 104782 65618 104866 65854
rect 105102 65618 105134 65854
rect 104514 26174 105134 65618
rect 104514 25938 104546 26174
rect 104782 25938 104866 26174
rect 105102 25938 105134 26174
rect 104514 25854 105134 25938
rect 104514 25618 104546 25854
rect 104782 25618 104866 25854
rect 105102 25618 105134 25854
rect 104514 -3226 105134 25618
rect 104514 -3462 104546 -3226
rect 104782 -3462 104866 -3226
rect 105102 -3462 105134 -3226
rect 104514 -3546 105134 -3462
rect 104514 -3782 104546 -3546
rect 104782 -3782 104866 -3546
rect 105102 -3782 105134 -3546
rect 104514 -3814 105134 -3782
rect 108234 669894 108854 709082
rect 108234 669658 108266 669894
rect 108502 669658 108586 669894
rect 108822 669658 108854 669894
rect 108234 669574 108854 669658
rect 108234 669338 108266 669574
rect 108502 669338 108586 669574
rect 108822 669338 108854 669574
rect 108234 629894 108854 669338
rect 108234 629658 108266 629894
rect 108502 629658 108586 629894
rect 108822 629658 108854 629894
rect 108234 629574 108854 629658
rect 108234 629338 108266 629574
rect 108502 629338 108586 629574
rect 108822 629338 108854 629574
rect 108234 589894 108854 629338
rect 108234 589658 108266 589894
rect 108502 589658 108586 589894
rect 108822 589658 108854 589894
rect 108234 589574 108854 589658
rect 108234 589338 108266 589574
rect 108502 589338 108586 589574
rect 108822 589338 108854 589574
rect 108234 549894 108854 589338
rect 108234 549658 108266 549894
rect 108502 549658 108586 549894
rect 108822 549658 108854 549894
rect 108234 549574 108854 549658
rect 108234 549338 108266 549574
rect 108502 549338 108586 549574
rect 108822 549338 108854 549574
rect 108234 509894 108854 549338
rect 108234 509658 108266 509894
rect 108502 509658 108586 509894
rect 108822 509658 108854 509894
rect 108234 509574 108854 509658
rect 108234 509338 108266 509574
rect 108502 509338 108586 509574
rect 108822 509338 108854 509574
rect 108234 469894 108854 509338
rect 108234 469658 108266 469894
rect 108502 469658 108586 469894
rect 108822 469658 108854 469894
rect 108234 469574 108854 469658
rect 108234 469338 108266 469574
rect 108502 469338 108586 469574
rect 108822 469338 108854 469574
rect 108234 429894 108854 469338
rect 108234 429658 108266 429894
rect 108502 429658 108586 429894
rect 108822 429658 108854 429894
rect 108234 429574 108854 429658
rect 108234 429338 108266 429574
rect 108502 429338 108586 429574
rect 108822 429338 108854 429574
rect 108234 389894 108854 429338
rect 108234 389658 108266 389894
rect 108502 389658 108586 389894
rect 108822 389658 108854 389894
rect 108234 389574 108854 389658
rect 108234 389338 108266 389574
rect 108502 389338 108586 389574
rect 108822 389338 108854 389574
rect 108234 349894 108854 389338
rect 108234 349658 108266 349894
rect 108502 349658 108586 349894
rect 108822 349658 108854 349894
rect 108234 349574 108854 349658
rect 108234 349338 108266 349574
rect 108502 349338 108586 349574
rect 108822 349338 108854 349574
rect 108234 309894 108854 349338
rect 108234 309658 108266 309894
rect 108502 309658 108586 309894
rect 108822 309658 108854 309894
rect 108234 309574 108854 309658
rect 108234 309338 108266 309574
rect 108502 309338 108586 309574
rect 108822 309338 108854 309574
rect 108234 269894 108854 309338
rect 108234 269658 108266 269894
rect 108502 269658 108586 269894
rect 108822 269658 108854 269894
rect 108234 269574 108854 269658
rect 108234 269338 108266 269574
rect 108502 269338 108586 269574
rect 108822 269338 108854 269574
rect 108234 229894 108854 269338
rect 108234 229658 108266 229894
rect 108502 229658 108586 229894
rect 108822 229658 108854 229894
rect 108234 229574 108854 229658
rect 108234 229338 108266 229574
rect 108502 229338 108586 229574
rect 108822 229338 108854 229574
rect 108234 189894 108854 229338
rect 108234 189658 108266 189894
rect 108502 189658 108586 189894
rect 108822 189658 108854 189894
rect 108234 189574 108854 189658
rect 108234 189338 108266 189574
rect 108502 189338 108586 189574
rect 108822 189338 108854 189574
rect 108234 149894 108854 189338
rect 108234 149658 108266 149894
rect 108502 149658 108586 149894
rect 108822 149658 108854 149894
rect 108234 149574 108854 149658
rect 108234 149338 108266 149574
rect 108502 149338 108586 149574
rect 108822 149338 108854 149574
rect 108234 109894 108854 149338
rect 108234 109658 108266 109894
rect 108502 109658 108586 109894
rect 108822 109658 108854 109894
rect 108234 109574 108854 109658
rect 108234 109338 108266 109574
rect 108502 109338 108586 109574
rect 108822 109338 108854 109574
rect 108234 69894 108854 109338
rect 108234 69658 108266 69894
rect 108502 69658 108586 69894
rect 108822 69658 108854 69894
rect 108234 69574 108854 69658
rect 108234 69338 108266 69574
rect 108502 69338 108586 69574
rect 108822 69338 108854 69574
rect 108234 29894 108854 69338
rect 108234 29658 108266 29894
rect 108502 29658 108586 29894
rect 108822 29658 108854 29894
rect 108234 29574 108854 29658
rect 108234 29338 108266 29574
rect 108502 29338 108586 29574
rect 108822 29338 108854 29574
rect 108234 -5146 108854 29338
rect 108234 -5382 108266 -5146
rect 108502 -5382 108586 -5146
rect 108822 -5382 108854 -5146
rect 108234 -5466 108854 -5382
rect 108234 -5702 108266 -5466
rect 108502 -5702 108586 -5466
rect 108822 -5702 108854 -5466
rect 108234 -5734 108854 -5702
rect 111954 673614 112574 711002
rect 131954 710598 132574 711590
rect 131954 710362 131986 710598
rect 132222 710362 132306 710598
rect 132542 710362 132574 710598
rect 131954 710278 132574 710362
rect 131954 710042 131986 710278
rect 132222 710042 132306 710278
rect 132542 710042 132574 710278
rect 128234 708678 128854 709670
rect 128234 708442 128266 708678
rect 128502 708442 128586 708678
rect 128822 708442 128854 708678
rect 128234 708358 128854 708442
rect 128234 708122 128266 708358
rect 128502 708122 128586 708358
rect 128822 708122 128854 708358
rect 124514 706758 125134 707750
rect 124514 706522 124546 706758
rect 124782 706522 124866 706758
rect 125102 706522 125134 706758
rect 124514 706438 125134 706522
rect 124514 706202 124546 706438
rect 124782 706202 124866 706438
rect 125102 706202 125134 706438
rect 111954 673378 111986 673614
rect 112222 673378 112306 673614
rect 112542 673378 112574 673614
rect 111954 673294 112574 673378
rect 111954 673058 111986 673294
rect 112222 673058 112306 673294
rect 112542 673058 112574 673294
rect 111954 633614 112574 673058
rect 111954 633378 111986 633614
rect 112222 633378 112306 633614
rect 112542 633378 112574 633614
rect 111954 633294 112574 633378
rect 111954 633058 111986 633294
rect 112222 633058 112306 633294
rect 112542 633058 112574 633294
rect 111954 593614 112574 633058
rect 111954 593378 111986 593614
rect 112222 593378 112306 593614
rect 112542 593378 112574 593614
rect 111954 593294 112574 593378
rect 111954 593058 111986 593294
rect 112222 593058 112306 593294
rect 112542 593058 112574 593294
rect 111954 553614 112574 593058
rect 111954 553378 111986 553614
rect 112222 553378 112306 553614
rect 112542 553378 112574 553614
rect 111954 553294 112574 553378
rect 111954 553058 111986 553294
rect 112222 553058 112306 553294
rect 112542 553058 112574 553294
rect 111954 513614 112574 553058
rect 111954 513378 111986 513614
rect 112222 513378 112306 513614
rect 112542 513378 112574 513614
rect 111954 513294 112574 513378
rect 111954 513058 111986 513294
rect 112222 513058 112306 513294
rect 112542 513058 112574 513294
rect 111954 473614 112574 513058
rect 111954 473378 111986 473614
rect 112222 473378 112306 473614
rect 112542 473378 112574 473614
rect 111954 473294 112574 473378
rect 111954 473058 111986 473294
rect 112222 473058 112306 473294
rect 112542 473058 112574 473294
rect 111954 433614 112574 473058
rect 111954 433378 111986 433614
rect 112222 433378 112306 433614
rect 112542 433378 112574 433614
rect 111954 433294 112574 433378
rect 111954 433058 111986 433294
rect 112222 433058 112306 433294
rect 112542 433058 112574 433294
rect 111954 393614 112574 433058
rect 111954 393378 111986 393614
rect 112222 393378 112306 393614
rect 112542 393378 112574 393614
rect 111954 393294 112574 393378
rect 111954 393058 111986 393294
rect 112222 393058 112306 393294
rect 112542 393058 112574 393294
rect 111954 353614 112574 393058
rect 111954 353378 111986 353614
rect 112222 353378 112306 353614
rect 112542 353378 112574 353614
rect 111954 353294 112574 353378
rect 111954 353058 111986 353294
rect 112222 353058 112306 353294
rect 112542 353058 112574 353294
rect 111954 313614 112574 353058
rect 111954 313378 111986 313614
rect 112222 313378 112306 313614
rect 112542 313378 112574 313614
rect 111954 313294 112574 313378
rect 111954 313058 111986 313294
rect 112222 313058 112306 313294
rect 112542 313058 112574 313294
rect 111954 273614 112574 313058
rect 111954 273378 111986 273614
rect 112222 273378 112306 273614
rect 112542 273378 112574 273614
rect 111954 273294 112574 273378
rect 111954 273058 111986 273294
rect 112222 273058 112306 273294
rect 112542 273058 112574 273294
rect 111954 233614 112574 273058
rect 111954 233378 111986 233614
rect 112222 233378 112306 233614
rect 112542 233378 112574 233614
rect 111954 233294 112574 233378
rect 111954 233058 111986 233294
rect 112222 233058 112306 233294
rect 112542 233058 112574 233294
rect 111954 193614 112574 233058
rect 111954 193378 111986 193614
rect 112222 193378 112306 193614
rect 112542 193378 112574 193614
rect 111954 193294 112574 193378
rect 111954 193058 111986 193294
rect 112222 193058 112306 193294
rect 112542 193058 112574 193294
rect 111954 153614 112574 193058
rect 111954 153378 111986 153614
rect 112222 153378 112306 153614
rect 112542 153378 112574 153614
rect 111954 153294 112574 153378
rect 111954 153058 111986 153294
rect 112222 153058 112306 153294
rect 112542 153058 112574 153294
rect 111954 113614 112574 153058
rect 111954 113378 111986 113614
rect 112222 113378 112306 113614
rect 112542 113378 112574 113614
rect 111954 113294 112574 113378
rect 111954 113058 111986 113294
rect 112222 113058 112306 113294
rect 112542 113058 112574 113294
rect 111954 73614 112574 113058
rect 111954 73378 111986 73614
rect 112222 73378 112306 73614
rect 112542 73378 112574 73614
rect 111954 73294 112574 73378
rect 111954 73058 111986 73294
rect 112222 73058 112306 73294
rect 112542 73058 112574 73294
rect 111954 33614 112574 73058
rect 111954 33378 111986 33614
rect 112222 33378 112306 33614
rect 112542 33378 112574 33614
rect 111954 33294 112574 33378
rect 111954 33058 111986 33294
rect 112222 33058 112306 33294
rect 112542 33058 112574 33294
rect 91954 -6342 91986 -6106
rect 92222 -6342 92306 -6106
rect 92542 -6342 92574 -6106
rect 91954 -6426 92574 -6342
rect 91954 -6662 91986 -6426
rect 92222 -6662 92306 -6426
rect 92542 -6662 92574 -6426
rect 91954 -7654 92574 -6662
rect 111954 -7066 112574 33058
rect 120794 704838 121414 705830
rect 120794 704602 120826 704838
rect 121062 704602 121146 704838
rect 121382 704602 121414 704838
rect 120794 704518 121414 704602
rect 120794 704282 120826 704518
rect 121062 704282 121146 704518
rect 121382 704282 121414 704518
rect 120794 682454 121414 704282
rect 120794 682218 120826 682454
rect 121062 682218 121146 682454
rect 121382 682218 121414 682454
rect 120794 682134 121414 682218
rect 120794 681898 120826 682134
rect 121062 681898 121146 682134
rect 121382 681898 121414 682134
rect 120794 642454 121414 681898
rect 120794 642218 120826 642454
rect 121062 642218 121146 642454
rect 121382 642218 121414 642454
rect 120794 642134 121414 642218
rect 120794 641898 120826 642134
rect 121062 641898 121146 642134
rect 121382 641898 121414 642134
rect 120794 602454 121414 641898
rect 120794 602218 120826 602454
rect 121062 602218 121146 602454
rect 121382 602218 121414 602454
rect 120794 602134 121414 602218
rect 120794 601898 120826 602134
rect 121062 601898 121146 602134
rect 121382 601898 121414 602134
rect 120794 562454 121414 601898
rect 120794 562218 120826 562454
rect 121062 562218 121146 562454
rect 121382 562218 121414 562454
rect 120794 562134 121414 562218
rect 120794 561898 120826 562134
rect 121062 561898 121146 562134
rect 121382 561898 121414 562134
rect 120794 522454 121414 561898
rect 120794 522218 120826 522454
rect 121062 522218 121146 522454
rect 121382 522218 121414 522454
rect 120794 522134 121414 522218
rect 120794 521898 120826 522134
rect 121062 521898 121146 522134
rect 121382 521898 121414 522134
rect 120794 482454 121414 521898
rect 120794 482218 120826 482454
rect 121062 482218 121146 482454
rect 121382 482218 121414 482454
rect 120794 482134 121414 482218
rect 120794 481898 120826 482134
rect 121062 481898 121146 482134
rect 121382 481898 121414 482134
rect 120794 442454 121414 481898
rect 120794 442218 120826 442454
rect 121062 442218 121146 442454
rect 121382 442218 121414 442454
rect 120794 442134 121414 442218
rect 120794 441898 120826 442134
rect 121062 441898 121146 442134
rect 121382 441898 121414 442134
rect 120794 402454 121414 441898
rect 120794 402218 120826 402454
rect 121062 402218 121146 402454
rect 121382 402218 121414 402454
rect 120794 402134 121414 402218
rect 120794 401898 120826 402134
rect 121062 401898 121146 402134
rect 121382 401898 121414 402134
rect 120794 362454 121414 401898
rect 120794 362218 120826 362454
rect 121062 362218 121146 362454
rect 121382 362218 121414 362454
rect 120794 362134 121414 362218
rect 120794 361898 120826 362134
rect 121062 361898 121146 362134
rect 121382 361898 121414 362134
rect 120794 322454 121414 361898
rect 120794 322218 120826 322454
rect 121062 322218 121146 322454
rect 121382 322218 121414 322454
rect 120794 322134 121414 322218
rect 120794 321898 120826 322134
rect 121062 321898 121146 322134
rect 121382 321898 121414 322134
rect 120794 282454 121414 321898
rect 120794 282218 120826 282454
rect 121062 282218 121146 282454
rect 121382 282218 121414 282454
rect 120794 282134 121414 282218
rect 120794 281898 120826 282134
rect 121062 281898 121146 282134
rect 121382 281898 121414 282134
rect 120794 242454 121414 281898
rect 120794 242218 120826 242454
rect 121062 242218 121146 242454
rect 121382 242218 121414 242454
rect 120794 242134 121414 242218
rect 120794 241898 120826 242134
rect 121062 241898 121146 242134
rect 121382 241898 121414 242134
rect 120794 202454 121414 241898
rect 120794 202218 120826 202454
rect 121062 202218 121146 202454
rect 121382 202218 121414 202454
rect 120794 202134 121414 202218
rect 120794 201898 120826 202134
rect 121062 201898 121146 202134
rect 121382 201898 121414 202134
rect 120794 162454 121414 201898
rect 120794 162218 120826 162454
rect 121062 162218 121146 162454
rect 121382 162218 121414 162454
rect 120794 162134 121414 162218
rect 120794 161898 120826 162134
rect 121062 161898 121146 162134
rect 121382 161898 121414 162134
rect 120794 122454 121414 161898
rect 120794 122218 120826 122454
rect 121062 122218 121146 122454
rect 121382 122218 121414 122454
rect 120794 122134 121414 122218
rect 120794 121898 120826 122134
rect 121062 121898 121146 122134
rect 121382 121898 121414 122134
rect 120794 82454 121414 121898
rect 120794 82218 120826 82454
rect 121062 82218 121146 82454
rect 121382 82218 121414 82454
rect 120794 82134 121414 82218
rect 120794 81898 120826 82134
rect 121062 81898 121146 82134
rect 121382 81898 121414 82134
rect 120794 42454 121414 81898
rect 120794 42218 120826 42454
rect 121062 42218 121146 42454
rect 121382 42218 121414 42454
rect 120794 42134 121414 42218
rect 120794 41898 120826 42134
rect 121062 41898 121146 42134
rect 121382 41898 121414 42134
rect 120794 2454 121414 41898
rect 120794 2218 120826 2454
rect 121062 2218 121146 2454
rect 121382 2218 121414 2454
rect 120794 2134 121414 2218
rect 120794 1898 120826 2134
rect 121062 1898 121146 2134
rect 121382 1898 121414 2134
rect 120794 -346 121414 1898
rect 120794 -582 120826 -346
rect 121062 -582 121146 -346
rect 121382 -582 121414 -346
rect 120794 -666 121414 -582
rect 120794 -902 120826 -666
rect 121062 -902 121146 -666
rect 121382 -902 121414 -666
rect 120794 -1894 121414 -902
rect 124514 686174 125134 706202
rect 124514 685938 124546 686174
rect 124782 685938 124866 686174
rect 125102 685938 125134 686174
rect 124514 685854 125134 685938
rect 124514 685618 124546 685854
rect 124782 685618 124866 685854
rect 125102 685618 125134 685854
rect 124514 646174 125134 685618
rect 124514 645938 124546 646174
rect 124782 645938 124866 646174
rect 125102 645938 125134 646174
rect 124514 645854 125134 645938
rect 124514 645618 124546 645854
rect 124782 645618 124866 645854
rect 125102 645618 125134 645854
rect 124514 606174 125134 645618
rect 124514 605938 124546 606174
rect 124782 605938 124866 606174
rect 125102 605938 125134 606174
rect 124514 605854 125134 605938
rect 124514 605618 124546 605854
rect 124782 605618 124866 605854
rect 125102 605618 125134 605854
rect 124514 566174 125134 605618
rect 124514 565938 124546 566174
rect 124782 565938 124866 566174
rect 125102 565938 125134 566174
rect 124514 565854 125134 565938
rect 124514 565618 124546 565854
rect 124782 565618 124866 565854
rect 125102 565618 125134 565854
rect 124514 526174 125134 565618
rect 124514 525938 124546 526174
rect 124782 525938 124866 526174
rect 125102 525938 125134 526174
rect 124514 525854 125134 525938
rect 124514 525618 124546 525854
rect 124782 525618 124866 525854
rect 125102 525618 125134 525854
rect 124514 486174 125134 525618
rect 124514 485938 124546 486174
rect 124782 485938 124866 486174
rect 125102 485938 125134 486174
rect 124514 485854 125134 485938
rect 124514 485618 124546 485854
rect 124782 485618 124866 485854
rect 125102 485618 125134 485854
rect 124514 446174 125134 485618
rect 124514 445938 124546 446174
rect 124782 445938 124866 446174
rect 125102 445938 125134 446174
rect 124514 445854 125134 445938
rect 124514 445618 124546 445854
rect 124782 445618 124866 445854
rect 125102 445618 125134 445854
rect 124514 406174 125134 445618
rect 124514 405938 124546 406174
rect 124782 405938 124866 406174
rect 125102 405938 125134 406174
rect 124514 405854 125134 405938
rect 124514 405618 124546 405854
rect 124782 405618 124866 405854
rect 125102 405618 125134 405854
rect 124514 366174 125134 405618
rect 124514 365938 124546 366174
rect 124782 365938 124866 366174
rect 125102 365938 125134 366174
rect 124514 365854 125134 365938
rect 124514 365618 124546 365854
rect 124782 365618 124866 365854
rect 125102 365618 125134 365854
rect 124514 326174 125134 365618
rect 124514 325938 124546 326174
rect 124782 325938 124866 326174
rect 125102 325938 125134 326174
rect 124514 325854 125134 325938
rect 124514 325618 124546 325854
rect 124782 325618 124866 325854
rect 125102 325618 125134 325854
rect 124514 286174 125134 325618
rect 124514 285938 124546 286174
rect 124782 285938 124866 286174
rect 125102 285938 125134 286174
rect 124514 285854 125134 285938
rect 124514 285618 124546 285854
rect 124782 285618 124866 285854
rect 125102 285618 125134 285854
rect 124514 246174 125134 285618
rect 124514 245938 124546 246174
rect 124782 245938 124866 246174
rect 125102 245938 125134 246174
rect 124514 245854 125134 245938
rect 124514 245618 124546 245854
rect 124782 245618 124866 245854
rect 125102 245618 125134 245854
rect 124514 206174 125134 245618
rect 124514 205938 124546 206174
rect 124782 205938 124866 206174
rect 125102 205938 125134 206174
rect 124514 205854 125134 205938
rect 124514 205618 124546 205854
rect 124782 205618 124866 205854
rect 125102 205618 125134 205854
rect 124514 166174 125134 205618
rect 124514 165938 124546 166174
rect 124782 165938 124866 166174
rect 125102 165938 125134 166174
rect 124514 165854 125134 165938
rect 124514 165618 124546 165854
rect 124782 165618 124866 165854
rect 125102 165618 125134 165854
rect 124514 126174 125134 165618
rect 124514 125938 124546 126174
rect 124782 125938 124866 126174
rect 125102 125938 125134 126174
rect 124514 125854 125134 125938
rect 124514 125618 124546 125854
rect 124782 125618 124866 125854
rect 125102 125618 125134 125854
rect 124514 86174 125134 125618
rect 124514 85938 124546 86174
rect 124782 85938 124866 86174
rect 125102 85938 125134 86174
rect 124514 85854 125134 85938
rect 124514 85618 124546 85854
rect 124782 85618 124866 85854
rect 125102 85618 125134 85854
rect 124514 46174 125134 85618
rect 124514 45938 124546 46174
rect 124782 45938 124866 46174
rect 125102 45938 125134 46174
rect 124514 45854 125134 45938
rect 124514 45618 124546 45854
rect 124782 45618 124866 45854
rect 125102 45618 125134 45854
rect 124514 6174 125134 45618
rect 124514 5938 124546 6174
rect 124782 5938 124866 6174
rect 125102 5938 125134 6174
rect 124514 5854 125134 5938
rect 124514 5618 124546 5854
rect 124782 5618 124866 5854
rect 125102 5618 125134 5854
rect 124514 -2266 125134 5618
rect 124514 -2502 124546 -2266
rect 124782 -2502 124866 -2266
rect 125102 -2502 125134 -2266
rect 124514 -2586 125134 -2502
rect 124514 -2822 124546 -2586
rect 124782 -2822 124866 -2586
rect 125102 -2822 125134 -2586
rect 124514 -3814 125134 -2822
rect 128234 689894 128854 708122
rect 128234 689658 128266 689894
rect 128502 689658 128586 689894
rect 128822 689658 128854 689894
rect 128234 689574 128854 689658
rect 128234 689338 128266 689574
rect 128502 689338 128586 689574
rect 128822 689338 128854 689574
rect 128234 649894 128854 689338
rect 128234 649658 128266 649894
rect 128502 649658 128586 649894
rect 128822 649658 128854 649894
rect 128234 649574 128854 649658
rect 128234 649338 128266 649574
rect 128502 649338 128586 649574
rect 128822 649338 128854 649574
rect 128234 609894 128854 649338
rect 128234 609658 128266 609894
rect 128502 609658 128586 609894
rect 128822 609658 128854 609894
rect 128234 609574 128854 609658
rect 128234 609338 128266 609574
rect 128502 609338 128586 609574
rect 128822 609338 128854 609574
rect 128234 569894 128854 609338
rect 128234 569658 128266 569894
rect 128502 569658 128586 569894
rect 128822 569658 128854 569894
rect 128234 569574 128854 569658
rect 128234 569338 128266 569574
rect 128502 569338 128586 569574
rect 128822 569338 128854 569574
rect 128234 529894 128854 569338
rect 128234 529658 128266 529894
rect 128502 529658 128586 529894
rect 128822 529658 128854 529894
rect 128234 529574 128854 529658
rect 128234 529338 128266 529574
rect 128502 529338 128586 529574
rect 128822 529338 128854 529574
rect 128234 489894 128854 529338
rect 128234 489658 128266 489894
rect 128502 489658 128586 489894
rect 128822 489658 128854 489894
rect 128234 489574 128854 489658
rect 128234 489338 128266 489574
rect 128502 489338 128586 489574
rect 128822 489338 128854 489574
rect 128234 449894 128854 489338
rect 128234 449658 128266 449894
rect 128502 449658 128586 449894
rect 128822 449658 128854 449894
rect 128234 449574 128854 449658
rect 128234 449338 128266 449574
rect 128502 449338 128586 449574
rect 128822 449338 128854 449574
rect 128234 409894 128854 449338
rect 128234 409658 128266 409894
rect 128502 409658 128586 409894
rect 128822 409658 128854 409894
rect 128234 409574 128854 409658
rect 128234 409338 128266 409574
rect 128502 409338 128586 409574
rect 128822 409338 128854 409574
rect 128234 369894 128854 409338
rect 128234 369658 128266 369894
rect 128502 369658 128586 369894
rect 128822 369658 128854 369894
rect 128234 369574 128854 369658
rect 128234 369338 128266 369574
rect 128502 369338 128586 369574
rect 128822 369338 128854 369574
rect 128234 329894 128854 369338
rect 128234 329658 128266 329894
rect 128502 329658 128586 329894
rect 128822 329658 128854 329894
rect 128234 329574 128854 329658
rect 128234 329338 128266 329574
rect 128502 329338 128586 329574
rect 128822 329338 128854 329574
rect 128234 289894 128854 329338
rect 128234 289658 128266 289894
rect 128502 289658 128586 289894
rect 128822 289658 128854 289894
rect 128234 289574 128854 289658
rect 128234 289338 128266 289574
rect 128502 289338 128586 289574
rect 128822 289338 128854 289574
rect 128234 249894 128854 289338
rect 128234 249658 128266 249894
rect 128502 249658 128586 249894
rect 128822 249658 128854 249894
rect 128234 249574 128854 249658
rect 128234 249338 128266 249574
rect 128502 249338 128586 249574
rect 128822 249338 128854 249574
rect 128234 209894 128854 249338
rect 128234 209658 128266 209894
rect 128502 209658 128586 209894
rect 128822 209658 128854 209894
rect 128234 209574 128854 209658
rect 128234 209338 128266 209574
rect 128502 209338 128586 209574
rect 128822 209338 128854 209574
rect 128234 169894 128854 209338
rect 128234 169658 128266 169894
rect 128502 169658 128586 169894
rect 128822 169658 128854 169894
rect 128234 169574 128854 169658
rect 128234 169338 128266 169574
rect 128502 169338 128586 169574
rect 128822 169338 128854 169574
rect 128234 129894 128854 169338
rect 128234 129658 128266 129894
rect 128502 129658 128586 129894
rect 128822 129658 128854 129894
rect 128234 129574 128854 129658
rect 128234 129338 128266 129574
rect 128502 129338 128586 129574
rect 128822 129338 128854 129574
rect 128234 89894 128854 129338
rect 128234 89658 128266 89894
rect 128502 89658 128586 89894
rect 128822 89658 128854 89894
rect 128234 89574 128854 89658
rect 128234 89338 128266 89574
rect 128502 89338 128586 89574
rect 128822 89338 128854 89574
rect 128234 49894 128854 89338
rect 128234 49658 128266 49894
rect 128502 49658 128586 49894
rect 128822 49658 128854 49894
rect 128234 49574 128854 49658
rect 128234 49338 128266 49574
rect 128502 49338 128586 49574
rect 128822 49338 128854 49574
rect 128234 9894 128854 49338
rect 128234 9658 128266 9894
rect 128502 9658 128586 9894
rect 128822 9658 128854 9894
rect 128234 9574 128854 9658
rect 128234 9338 128266 9574
rect 128502 9338 128586 9574
rect 128822 9338 128854 9574
rect 128234 -4186 128854 9338
rect 128234 -4422 128266 -4186
rect 128502 -4422 128586 -4186
rect 128822 -4422 128854 -4186
rect 128234 -4506 128854 -4422
rect 128234 -4742 128266 -4506
rect 128502 -4742 128586 -4506
rect 128822 -4742 128854 -4506
rect 128234 -5734 128854 -4742
rect 131954 693614 132574 710042
rect 151954 711558 152574 711590
rect 151954 711322 151986 711558
rect 152222 711322 152306 711558
rect 152542 711322 152574 711558
rect 151954 711238 152574 711322
rect 151954 711002 151986 711238
rect 152222 711002 152306 711238
rect 152542 711002 152574 711238
rect 148234 709638 148854 709670
rect 148234 709402 148266 709638
rect 148502 709402 148586 709638
rect 148822 709402 148854 709638
rect 148234 709318 148854 709402
rect 148234 709082 148266 709318
rect 148502 709082 148586 709318
rect 148822 709082 148854 709318
rect 144514 707718 145134 707750
rect 144514 707482 144546 707718
rect 144782 707482 144866 707718
rect 145102 707482 145134 707718
rect 144514 707398 145134 707482
rect 144514 707162 144546 707398
rect 144782 707162 144866 707398
rect 145102 707162 145134 707398
rect 131954 693378 131986 693614
rect 132222 693378 132306 693614
rect 132542 693378 132574 693614
rect 131954 693294 132574 693378
rect 131954 693058 131986 693294
rect 132222 693058 132306 693294
rect 132542 693058 132574 693294
rect 131954 653614 132574 693058
rect 131954 653378 131986 653614
rect 132222 653378 132306 653614
rect 132542 653378 132574 653614
rect 131954 653294 132574 653378
rect 131954 653058 131986 653294
rect 132222 653058 132306 653294
rect 132542 653058 132574 653294
rect 131954 613614 132574 653058
rect 131954 613378 131986 613614
rect 132222 613378 132306 613614
rect 132542 613378 132574 613614
rect 131954 613294 132574 613378
rect 131954 613058 131986 613294
rect 132222 613058 132306 613294
rect 132542 613058 132574 613294
rect 131954 573614 132574 613058
rect 131954 573378 131986 573614
rect 132222 573378 132306 573614
rect 132542 573378 132574 573614
rect 131954 573294 132574 573378
rect 131954 573058 131986 573294
rect 132222 573058 132306 573294
rect 132542 573058 132574 573294
rect 131954 533614 132574 573058
rect 131954 533378 131986 533614
rect 132222 533378 132306 533614
rect 132542 533378 132574 533614
rect 131954 533294 132574 533378
rect 131954 533058 131986 533294
rect 132222 533058 132306 533294
rect 132542 533058 132574 533294
rect 131954 493614 132574 533058
rect 131954 493378 131986 493614
rect 132222 493378 132306 493614
rect 132542 493378 132574 493614
rect 131954 493294 132574 493378
rect 131954 493058 131986 493294
rect 132222 493058 132306 493294
rect 132542 493058 132574 493294
rect 131954 453614 132574 493058
rect 131954 453378 131986 453614
rect 132222 453378 132306 453614
rect 132542 453378 132574 453614
rect 131954 453294 132574 453378
rect 131954 453058 131986 453294
rect 132222 453058 132306 453294
rect 132542 453058 132574 453294
rect 131954 413614 132574 453058
rect 131954 413378 131986 413614
rect 132222 413378 132306 413614
rect 132542 413378 132574 413614
rect 131954 413294 132574 413378
rect 131954 413058 131986 413294
rect 132222 413058 132306 413294
rect 132542 413058 132574 413294
rect 131954 373614 132574 413058
rect 131954 373378 131986 373614
rect 132222 373378 132306 373614
rect 132542 373378 132574 373614
rect 131954 373294 132574 373378
rect 131954 373058 131986 373294
rect 132222 373058 132306 373294
rect 132542 373058 132574 373294
rect 131954 333614 132574 373058
rect 131954 333378 131986 333614
rect 132222 333378 132306 333614
rect 132542 333378 132574 333614
rect 131954 333294 132574 333378
rect 131954 333058 131986 333294
rect 132222 333058 132306 333294
rect 132542 333058 132574 333294
rect 131954 293614 132574 333058
rect 140794 705798 141414 705830
rect 140794 705562 140826 705798
rect 141062 705562 141146 705798
rect 141382 705562 141414 705798
rect 140794 705478 141414 705562
rect 140794 705242 140826 705478
rect 141062 705242 141146 705478
rect 141382 705242 141414 705478
rect 140794 662454 141414 705242
rect 140794 662218 140826 662454
rect 141062 662218 141146 662454
rect 141382 662218 141414 662454
rect 140794 662134 141414 662218
rect 140794 661898 140826 662134
rect 141062 661898 141146 662134
rect 141382 661898 141414 662134
rect 140794 622454 141414 661898
rect 140794 622218 140826 622454
rect 141062 622218 141146 622454
rect 141382 622218 141414 622454
rect 140794 622134 141414 622218
rect 140794 621898 140826 622134
rect 141062 621898 141146 622134
rect 141382 621898 141414 622134
rect 140794 582454 141414 621898
rect 140794 582218 140826 582454
rect 141062 582218 141146 582454
rect 141382 582218 141414 582454
rect 140794 582134 141414 582218
rect 140794 581898 140826 582134
rect 141062 581898 141146 582134
rect 141382 581898 141414 582134
rect 140794 542454 141414 581898
rect 140794 542218 140826 542454
rect 141062 542218 141146 542454
rect 141382 542218 141414 542454
rect 140794 542134 141414 542218
rect 140794 541898 140826 542134
rect 141062 541898 141146 542134
rect 141382 541898 141414 542134
rect 140794 502454 141414 541898
rect 140794 502218 140826 502454
rect 141062 502218 141146 502454
rect 141382 502218 141414 502454
rect 140794 502134 141414 502218
rect 140794 501898 140826 502134
rect 141062 501898 141146 502134
rect 141382 501898 141414 502134
rect 140794 462454 141414 501898
rect 140794 462218 140826 462454
rect 141062 462218 141146 462454
rect 141382 462218 141414 462454
rect 140794 462134 141414 462218
rect 140794 461898 140826 462134
rect 141062 461898 141146 462134
rect 141382 461898 141414 462134
rect 140794 422454 141414 461898
rect 140794 422218 140826 422454
rect 141062 422218 141146 422454
rect 141382 422218 141414 422454
rect 140794 422134 141414 422218
rect 140794 421898 140826 422134
rect 141062 421898 141146 422134
rect 141382 421898 141414 422134
rect 140794 382454 141414 421898
rect 140794 382218 140826 382454
rect 141062 382218 141146 382454
rect 141382 382218 141414 382454
rect 140794 382134 141414 382218
rect 140794 381898 140826 382134
rect 141062 381898 141146 382134
rect 141382 381898 141414 382134
rect 140794 342454 141414 381898
rect 140794 342218 140826 342454
rect 141062 342218 141146 342454
rect 141382 342218 141414 342454
rect 140794 342134 141414 342218
rect 140794 341898 140826 342134
rect 141062 341898 141146 342134
rect 141382 341898 141414 342134
rect 139163 319428 139229 319429
rect 139163 319364 139164 319428
rect 139228 319364 139229 319428
rect 139163 319363 139229 319364
rect 131954 293378 131986 293614
rect 132222 293378 132306 293614
rect 132542 293378 132574 293614
rect 131954 293294 132574 293378
rect 131954 293058 131986 293294
rect 132222 293058 132306 293294
rect 132542 293058 132574 293294
rect 131954 253614 132574 293058
rect 131954 253378 131986 253614
rect 132222 253378 132306 253614
rect 132542 253378 132574 253614
rect 131954 253294 132574 253378
rect 131954 253058 131986 253294
rect 132222 253058 132306 253294
rect 132542 253058 132574 253294
rect 131954 213614 132574 253058
rect 131954 213378 131986 213614
rect 132222 213378 132306 213614
rect 132542 213378 132574 213614
rect 131954 213294 132574 213378
rect 131954 213058 131986 213294
rect 132222 213058 132306 213294
rect 132542 213058 132574 213294
rect 131954 173614 132574 213058
rect 131954 173378 131986 173614
rect 132222 173378 132306 173614
rect 132542 173378 132574 173614
rect 131954 173294 132574 173378
rect 131954 173058 131986 173294
rect 132222 173058 132306 173294
rect 132542 173058 132574 173294
rect 131954 133614 132574 173058
rect 131954 133378 131986 133614
rect 132222 133378 132306 133614
rect 132542 133378 132574 133614
rect 131954 133294 132574 133378
rect 131954 133058 131986 133294
rect 132222 133058 132306 133294
rect 132542 133058 132574 133294
rect 131954 93614 132574 133058
rect 131954 93378 131986 93614
rect 132222 93378 132306 93614
rect 132542 93378 132574 93614
rect 131954 93294 132574 93378
rect 131954 93058 131986 93294
rect 132222 93058 132306 93294
rect 132542 93058 132574 93294
rect 131954 53614 132574 93058
rect 131954 53378 131986 53614
rect 132222 53378 132306 53614
rect 132542 53378 132574 53614
rect 131954 53294 132574 53378
rect 131954 53058 131986 53294
rect 132222 53058 132306 53294
rect 132542 53058 132574 53294
rect 131954 13614 132574 53058
rect 131954 13378 131986 13614
rect 132222 13378 132306 13614
rect 132542 13378 132574 13614
rect 131954 13294 132574 13378
rect 131954 13058 131986 13294
rect 132222 13058 132306 13294
rect 132542 13058 132574 13294
rect 111954 -7302 111986 -7066
rect 112222 -7302 112306 -7066
rect 112542 -7302 112574 -7066
rect 111954 -7386 112574 -7302
rect 111954 -7622 111986 -7386
rect 112222 -7622 112306 -7386
rect 112542 -7622 112574 -7386
rect 111954 -7654 112574 -7622
rect 131954 -6106 132574 13058
rect 139166 3501 139226 319363
rect 140794 302454 141414 341898
rect 140794 302218 140826 302454
rect 141382 302218 141414 302454
rect 140794 302134 141414 302218
rect 140794 301898 140826 302134
rect 141382 301898 141414 302134
rect 140794 262454 141414 301898
rect 140794 262218 140826 262454
rect 141382 262218 141414 262454
rect 140794 262134 141414 262218
rect 140794 261898 140826 262134
rect 141382 261898 141414 262134
rect 140794 222454 141414 261898
rect 140794 222218 140826 222454
rect 141382 222218 141414 222454
rect 140794 222134 141414 222218
rect 140794 221898 140826 222134
rect 141382 221898 141414 222134
rect 140794 182454 141414 221898
rect 140794 182218 140826 182454
rect 141382 182218 141414 182454
rect 140794 182134 141414 182218
rect 140794 181898 140826 182134
rect 141382 181898 141414 182134
rect 140794 142454 141414 181898
rect 140794 142218 140826 142454
rect 141382 142218 141414 142454
rect 140794 142134 141414 142218
rect 140794 141898 140826 142134
rect 141382 141898 141414 142134
rect 140794 102454 141414 141898
rect 140794 102218 140826 102454
rect 141062 102218 141146 102454
rect 141382 102218 141414 102454
rect 140794 102134 141414 102218
rect 140794 101898 140826 102134
rect 141062 101898 141146 102134
rect 141382 101898 141414 102134
rect 140794 62454 141414 101898
rect 140794 62218 140826 62454
rect 141062 62218 141146 62454
rect 141382 62218 141414 62454
rect 140794 62134 141414 62218
rect 140794 61898 140826 62134
rect 141062 61898 141146 62134
rect 141382 61898 141414 62134
rect 140794 22454 141414 61898
rect 140794 22218 140826 22454
rect 141062 22218 141146 22454
rect 141382 22218 141414 22454
rect 140794 22134 141414 22218
rect 140794 21898 140826 22134
rect 141062 21898 141146 22134
rect 141382 21898 141414 22134
rect 139163 3500 139229 3501
rect 139163 3436 139164 3500
rect 139228 3436 139229 3500
rect 139163 3435 139229 3436
rect 140794 -1306 141414 21898
rect 140794 -1542 140826 -1306
rect 141062 -1542 141146 -1306
rect 141382 -1542 141414 -1306
rect 140794 -1626 141414 -1542
rect 140794 -1862 140826 -1626
rect 141062 -1862 141146 -1626
rect 141382 -1862 141414 -1626
rect 140794 -1894 141414 -1862
rect 144514 666174 145134 707162
rect 144514 665938 144546 666174
rect 144782 665938 144866 666174
rect 145102 665938 145134 666174
rect 144514 665854 145134 665938
rect 144514 665618 144546 665854
rect 144782 665618 144866 665854
rect 145102 665618 145134 665854
rect 144514 626174 145134 665618
rect 144514 625938 144546 626174
rect 144782 625938 144866 626174
rect 145102 625938 145134 626174
rect 144514 625854 145134 625938
rect 144514 625618 144546 625854
rect 144782 625618 144866 625854
rect 145102 625618 145134 625854
rect 144514 586174 145134 625618
rect 144514 585938 144546 586174
rect 144782 585938 144866 586174
rect 145102 585938 145134 586174
rect 144514 585854 145134 585938
rect 144514 585618 144546 585854
rect 144782 585618 144866 585854
rect 145102 585618 145134 585854
rect 144514 546174 145134 585618
rect 144514 545938 144546 546174
rect 144782 545938 144866 546174
rect 145102 545938 145134 546174
rect 144514 545854 145134 545938
rect 144514 545618 144546 545854
rect 144782 545618 144866 545854
rect 145102 545618 145134 545854
rect 144514 506174 145134 545618
rect 144514 505938 144546 506174
rect 144782 505938 144866 506174
rect 145102 505938 145134 506174
rect 144514 505854 145134 505938
rect 144514 505618 144546 505854
rect 144782 505618 144866 505854
rect 145102 505618 145134 505854
rect 144514 466174 145134 505618
rect 144514 465938 144546 466174
rect 144782 465938 144866 466174
rect 145102 465938 145134 466174
rect 144514 465854 145134 465938
rect 144514 465618 144546 465854
rect 144782 465618 144866 465854
rect 145102 465618 145134 465854
rect 144514 426174 145134 465618
rect 144514 425938 144546 426174
rect 144782 425938 144866 426174
rect 145102 425938 145134 426174
rect 144514 425854 145134 425938
rect 144514 425618 144546 425854
rect 144782 425618 144866 425854
rect 145102 425618 145134 425854
rect 144514 386174 145134 425618
rect 144514 385938 144546 386174
rect 144782 385938 144866 386174
rect 145102 385938 145134 386174
rect 144514 385854 145134 385938
rect 144514 385618 144546 385854
rect 144782 385618 144866 385854
rect 145102 385618 145134 385854
rect 144514 346174 145134 385618
rect 144514 345938 144546 346174
rect 144782 345938 144866 346174
rect 145102 345938 145134 346174
rect 144514 345854 145134 345938
rect 144514 345618 144546 345854
rect 144782 345618 144866 345854
rect 145102 345618 145134 345854
rect 144514 306174 145134 345618
rect 144514 305938 144546 306174
rect 144782 305938 144866 306174
rect 145102 305938 145134 306174
rect 144514 305854 145134 305938
rect 144514 305618 144546 305854
rect 144782 305618 144866 305854
rect 145102 305618 145134 305854
rect 144514 266174 145134 305618
rect 144514 265938 144546 266174
rect 144782 265938 144866 266174
rect 145102 265938 145134 266174
rect 144514 265854 145134 265938
rect 144514 265618 144546 265854
rect 144782 265618 144866 265854
rect 145102 265618 145134 265854
rect 144514 226174 145134 265618
rect 144514 225938 144546 226174
rect 144782 225938 144866 226174
rect 145102 225938 145134 226174
rect 144514 225854 145134 225938
rect 144514 225618 144546 225854
rect 144782 225618 144866 225854
rect 145102 225618 145134 225854
rect 144514 186174 145134 225618
rect 144514 185938 144546 186174
rect 144782 185938 144866 186174
rect 145102 185938 145134 186174
rect 144514 185854 145134 185938
rect 144514 185618 144546 185854
rect 144782 185618 144866 185854
rect 145102 185618 145134 185854
rect 144514 146174 145134 185618
rect 144514 145938 144546 146174
rect 144782 145938 144866 146174
rect 145102 145938 145134 146174
rect 144514 145854 145134 145938
rect 144514 145618 144546 145854
rect 144782 145618 144866 145854
rect 145102 145618 145134 145854
rect 144514 106174 145134 145618
rect 144514 105938 144546 106174
rect 144782 105938 144866 106174
rect 145102 105938 145134 106174
rect 144514 105854 145134 105938
rect 144514 105618 144546 105854
rect 144782 105618 144866 105854
rect 145102 105618 145134 105854
rect 144514 66174 145134 105618
rect 144514 65938 144546 66174
rect 144782 65938 144866 66174
rect 145102 65938 145134 66174
rect 144514 65854 145134 65938
rect 144514 65618 144546 65854
rect 144782 65618 144866 65854
rect 145102 65618 145134 65854
rect 144514 26174 145134 65618
rect 144514 25938 144546 26174
rect 144782 25938 144866 26174
rect 145102 25938 145134 26174
rect 144514 25854 145134 25938
rect 144514 25618 144546 25854
rect 144782 25618 144866 25854
rect 145102 25618 145134 25854
rect 144514 -3226 145134 25618
rect 144514 -3462 144546 -3226
rect 144782 -3462 144866 -3226
rect 145102 -3462 145134 -3226
rect 144514 -3546 145134 -3462
rect 144514 -3782 144546 -3546
rect 144782 -3782 144866 -3546
rect 145102 -3782 145134 -3546
rect 144514 -3814 145134 -3782
rect 148234 669894 148854 709082
rect 148234 669658 148266 669894
rect 148502 669658 148586 669894
rect 148822 669658 148854 669894
rect 148234 669574 148854 669658
rect 148234 669338 148266 669574
rect 148502 669338 148586 669574
rect 148822 669338 148854 669574
rect 148234 629894 148854 669338
rect 148234 629658 148266 629894
rect 148502 629658 148586 629894
rect 148822 629658 148854 629894
rect 148234 629574 148854 629658
rect 148234 629338 148266 629574
rect 148502 629338 148586 629574
rect 148822 629338 148854 629574
rect 148234 589894 148854 629338
rect 148234 589658 148266 589894
rect 148502 589658 148586 589894
rect 148822 589658 148854 589894
rect 148234 589574 148854 589658
rect 148234 589338 148266 589574
rect 148502 589338 148586 589574
rect 148822 589338 148854 589574
rect 148234 549894 148854 589338
rect 148234 549658 148266 549894
rect 148502 549658 148586 549894
rect 148822 549658 148854 549894
rect 148234 549574 148854 549658
rect 148234 549338 148266 549574
rect 148502 549338 148586 549574
rect 148822 549338 148854 549574
rect 148234 509894 148854 549338
rect 148234 509658 148266 509894
rect 148502 509658 148586 509894
rect 148822 509658 148854 509894
rect 148234 509574 148854 509658
rect 148234 509338 148266 509574
rect 148502 509338 148586 509574
rect 148822 509338 148854 509574
rect 148234 469894 148854 509338
rect 148234 469658 148266 469894
rect 148502 469658 148586 469894
rect 148822 469658 148854 469894
rect 148234 469574 148854 469658
rect 148234 469338 148266 469574
rect 148502 469338 148586 469574
rect 148822 469338 148854 469574
rect 148234 429894 148854 469338
rect 148234 429658 148266 429894
rect 148502 429658 148586 429894
rect 148822 429658 148854 429894
rect 148234 429574 148854 429658
rect 148234 429338 148266 429574
rect 148502 429338 148586 429574
rect 148822 429338 148854 429574
rect 148234 389894 148854 429338
rect 148234 389658 148266 389894
rect 148502 389658 148586 389894
rect 148822 389658 148854 389894
rect 148234 389574 148854 389658
rect 148234 389338 148266 389574
rect 148502 389338 148586 389574
rect 148822 389338 148854 389574
rect 148234 349894 148854 389338
rect 148234 349658 148266 349894
rect 148502 349658 148586 349894
rect 148822 349658 148854 349894
rect 148234 349574 148854 349658
rect 148234 349338 148266 349574
rect 148502 349338 148586 349574
rect 148822 349338 148854 349574
rect 148234 309894 148854 349338
rect 148234 309658 148266 309894
rect 148502 309658 148586 309894
rect 148822 309658 148854 309894
rect 148234 309574 148854 309658
rect 148234 309338 148266 309574
rect 148502 309338 148586 309574
rect 148822 309338 148854 309574
rect 148234 269894 148854 309338
rect 148234 269658 148266 269894
rect 148502 269658 148586 269894
rect 148822 269658 148854 269894
rect 148234 269574 148854 269658
rect 148234 269338 148266 269574
rect 148502 269338 148586 269574
rect 148822 269338 148854 269574
rect 148234 229894 148854 269338
rect 148234 229658 148266 229894
rect 148502 229658 148586 229894
rect 148822 229658 148854 229894
rect 148234 229574 148854 229658
rect 148234 229338 148266 229574
rect 148502 229338 148586 229574
rect 148822 229338 148854 229574
rect 148234 189894 148854 229338
rect 148234 189658 148266 189894
rect 148502 189658 148586 189894
rect 148822 189658 148854 189894
rect 148234 189574 148854 189658
rect 148234 189338 148266 189574
rect 148502 189338 148586 189574
rect 148822 189338 148854 189574
rect 148234 149894 148854 189338
rect 148234 149658 148266 149894
rect 148502 149658 148586 149894
rect 148822 149658 148854 149894
rect 148234 149574 148854 149658
rect 148234 149338 148266 149574
rect 148502 149338 148586 149574
rect 148822 149338 148854 149574
rect 148234 109894 148854 149338
rect 148234 109658 148266 109894
rect 148502 109658 148586 109894
rect 148822 109658 148854 109894
rect 148234 109574 148854 109658
rect 148234 109338 148266 109574
rect 148502 109338 148586 109574
rect 148822 109338 148854 109574
rect 148234 69894 148854 109338
rect 148234 69658 148266 69894
rect 148502 69658 148586 69894
rect 148822 69658 148854 69894
rect 148234 69574 148854 69658
rect 148234 69338 148266 69574
rect 148502 69338 148586 69574
rect 148822 69338 148854 69574
rect 148234 29894 148854 69338
rect 148234 29658 148266 29894
rect 148502 29658 148586 29894
rect 148822 29658 148854 29894
rect 148234 29574 148854 29658
rect 148234 29338 148266 29574
rect 148502 29338 148586 29574
rect 148822 29338 148854 29574
rect 148234 -5146 148854 29338
rect 148234 -5382 148266 -5146
rect 148502 -5382 148586 -5146
rect 148822 -5382 148854 -5146
rect 148234 -5466 148854 -5382
rect 148234 -5702 148266 -5466
rect 148502 -5702 148586 -5466
rect 148822 -5702 148854 -5466
rect 148234 -5734 148854 -5702
rect 151954 673614 152574 711002
rect 171954 710598 172574 711590
rect 171954 710362 171986 710598
rect 172222 710362 172306 710598
rect 172542 710362 172574 710598
rect 171954 710278 172574 710362
rect 171954 710042 171986 710278
rect 172222 710042 172306 710278
rect 172542 710042 172574 710278
rect 168234 708678 168854 709670
rect 168234 708442 168266 708678
rect 168502 708442 168586 708678
rect 168822 708442 168854 708678
rect 168234 708358 168854 708442
rect 168234 708122 168266 708358
rect 168502 708122 168586 708358
rect 168822 708122 168854 708358
rect 164514 706758 165134 707750
rect 164514 706522 164546 706758
rect 164782 706522 164866 706758
rect 165102 706522 165134 706758
rect 164514 706438 165134 706522
rect 164514 706202 164546 706438
rect 164782 706202 164866 706438
rect 165102 706202 165134 706438
rect 151954 673378 151986 673614
rect 152222 673378 152306 673614
rect 152542 673378 152574 673614
rect 151954 673294 152574 673378
rect 151954 673058 151986 673294
rect 152222 673058 152306 673294
rect 152542 673058 152574 673294
rect 151954 633614 152574 673058
rect 151954 633378 151986 633614
rect 152222 633378 152306 633614
rect 152542 633378 152574 633614
rect 151954 633294 152574 633378
rect 151954 633058 151986 633294
rect 152222 633058 152306 633294
rect 152542 633058 152574 633294
rect 151954 593614 152574 633058
rect 151954 593378 151986 593614
rect 152222 593378 152306 593614
rect 152542 593378 152574 593614
rect 151954 593294 152574 593378
rect 151954 593058 151986 593294
rect 152222 593058 152306 593294
rect 152542 593058 152574 593294
rect 151954 553614 152574 593058
rect 151954 553378 151986 553614
rect 152222 553378 152306 553614
rect 152542 553378 152574 553614
rect 151954 553294 152574 553378
rect 151954 553058 151986 553294
rect 152222 553058 152306 553294
rect 152542 553058 152574 553294
rect 151954 513614 152574 553058
rect 151954 513378 151986 513614
rect 152222 513378 152306 513614
rect 152542 513378 152574 513614
rect 151954 513294 152574 513378
rect 151954 513058 151986 513294
rect 152222 513058 152306 513294
rect 152542 513058 152574 513294
rect 151954 473614 152574 513058
rect 151954 473378 151986 473614
rect 152222 473378 152306 473614
rect 152542 473378 152574 473614
rect 151954 473294 152574 473378
rect 151954 473058 151986 473294
rect 152222 473058 152306 473294
rect 152542 473058 152574 473294
rect 151954 433614 152574 473058
rect 151954 433378 151986 433614
rect 152222 433378 152306 433614
rect 152542 433378 152574 433614
rect 151954 433294 152574 433378
rect 151954 433058 151986 433294
rect 152222 433058 152306 433294
rect 152542 433058 152574 433294
rect 151954 393614 152574 433058
rect 151954 393378 151986 393614
rect 152222 393378 152306 393614
rect 152542 393378 152574 393614
rect 151954 393294 152574 393378
rect 151954 393058 151986 393294
rect 152222 393058 152306 393294
rect 152542 393058 152574 393294
rect 151954 353614 152574 393058
rect 151954 353378 151986 353614
rect 152222 353378 152306 353614
rect 152542 353378 152574 353614
rect 151954 353294 152574 353378
rect 151954 353058 151986 353294
rect 152222 353058 152306 353294
rect 152542 353058 152574 353294
rect 151954 313614 152574 353058
rect 160794 704838 161414 705830
rect 160794 704602 160826 704838
rect 161062 704602 161146 704838
rect 161382 704602 161414 704838
rect 160794 704518 161414 704602
rect 160794 704282 160826 704518
rect 161062 704282 161146 704518
rect 161382 704282 161414 704518
rect 160794 682454 161414 704282
rect 160794 682218 160826 682454
rect 161062 682218 161146 682454
rect 161382 682218 161414 682454
rect 160794 682134 161414 682218
rect 160794 681898 160826 682134
rect 161062 681898 161146 682134
rect 161382 681898 161414 682134
rect 160794 642454 161414 681898
rect 160794 642218 160826 642454
rect 161062 642218 161146 642454
rect 161382 642218 161414 642454
rect 160794 642134 161414 642218
rect 160794 641898 160826 642134
rect 161062 641898 161146 642134
rect 161382 641898 161414 642134
rect 160794 602454 161414 641898
rect 160794 602218 160826 602454
rect 161062 602218 161146 602454
rect 161382 602218 161414 602454
rect 160794 602134 161414 602218
rect 160794 601898 160826 602134
rect 161062 601898 161146 602134
rect 161382 601898 161414 602134
rect 160794 562454 161414 601898
rect 160794 562218 160826 562454
rect 161062 562218 161146 562454
rect 161382 562218 161414 562454
rect 160794 562134 161414 562218
rect 160794 561898 160826 562134
rect 161062 561898 161146 562134
rect 161382 561898 161414 562134
rect 160794 522454 161414 561898
rect 160794 522218 160826 522454
rect 161062 522218 161146 522454
rect 161382 522218 161414 522454
rect 160794 522134 161414 522218
rect 160794 521898 160826 522134
rect 161062 521898 161146 522134
rect 161382 521898 161414 522134
rect 160794 482454 161414 521898
rect 160794 482218 160826 482454
rect 161062 482218 161146 482454
rect 161382 482218 161414 482454
rect 160794 482134 161414 482218
rect 160794 481898 160826 482134
rect 161062 481898 161146 482134
rect 161382 481898 161414 482134
rect 160794 442454 161414 481898
rect 160794 442218 160826 442454
rect 161062 442218 161146 442454
rect 161382 442218 161414 442454
rect 160794 442134 161414 442218
rect 160794 441898 160826 442134
rect 161062 441898 161146 442134
rect 161382 441898 161414 442134
rect 160794 402454 161414 441898
rect 160794 402218 160826 402454
rect 161062 402218 161146 402454
rect 161382 402218 161414 402454
rect 160794 402134 161414 402218
rect 160794 401898 160826 402134
rect 161062 401898 161146 402134
rect 161382 401898 161414 402134
rect 160794 362454 161414 401898
rect 160794 362218 160826 362454
rect 161062 362218 161146 362454
rect 161382 362218 161414 362454
rect 160794 362134 161414 362218
rect 160794 361898 160826 362134
rect 161062 361898 161146 362134
rect 161382 361898 161414 362134
rect 160794 322454 161414 361898
rect 160794 322218 160826 322454
rect 161062 322218 161146 322454
rect 161382 322218 161414 322454
rect 160794 322134 161414 322218
rect 160794 321898 160826 322134
rect 161062 321898 161146 322134
rect 161382 321898 161414 322134
rect 160507 319428 160573 319429
rect 160507 319364 160508 319428
rect 160572 319364 160573 319428
rect 160507 319363 160573 319364
rect 151954 313378 151986 313614
rect 152222 313378 152306 313614
rect 152542 313378 152574 313614
rect 151954 313294 152574 313378
rect 151954 313058 151986 313294
rect 152222 313058 152306 313294
rect 152542 313058 152574 313294
rect 151954 273614 152574 313058
rect 151954 273378 151986 273614
rect 152222 273378 152306 273614
rect 152542 273378 152574 273614
rect 151954 273294 152574 273378
rect 151954 273058 151986 273294
rect 152222 273058 152306 273294
rect 152542 273058 152574 273294
rect 151954 233614 152574 273058
rect 151954 233378 151986 233614
rect 152222 233378 152306 233614
rect 152542 233378 152574 233614
rect 151954 233294 152574 233378
rect 151954 233058 151986 233294
rect 152222 233058 152306 233294
rect 152542 233058 152574 233294
rect 151954 193614 152574 233058
rect 151954 193378 151986 193614
rect 152222 193378 152306 193614
rect 152542 193378 152574 193614
rect 151954 193294 152574 193378
rect 151954 193058 151986 193294
rect 152222 193058 152306 193294
rect 152542 193058 152574 193294
rect 151954 153614 152574 193058
rect 151954 153378 151986 153614
rect 152222 153378 152306 153614
rect 152542 153378 152574 153614
rect 151954 153294 152574 153378
rect 151954 153058 151986 153294
rect 152222 153058 152306 153294
rect 152542 153058 152574 153294
rect 151954 113614 152574 153058
rect 151954 113378 151986 113614
rect 152222 113378 152306 113614
rect 152542 113378 152574 113614
rect 151954 113294 152574 113378
rect 151954 113058 151986 113294
rect 152222 113058 152306 113294
rect 152542 113058 152574 113294
rect 151954 73614 152574 113058
rect 151954 73378 151986 73614
rect 152222 73378 152306 73614
rect 152542 73378 152574 73614
rect 151954 73294 152574 73378
rect 151954 73058 151986 73294
rect 152222 73058 152306 73294
rect 152542 73058 152574 73294
rect 151954 33614 152574 73058
rect 151954 33378 151986 33614
rect 152222 33378 152306 33614
rect 152542 33378 152574 33614
rect 151954 33294 152574 33378
rect 151954 33058 151986 33294
rect 152222 33058 152306 33294
rect 152542 33058 152574 33294
rect 131954 -6342 131986 -6106
rect 132222 -6342 132306 -6106
rect 132542 -6342 132574 -6106
rect 131954 -6426 132574 -6342
rect 131954 -6662 131986 -6426
rect 132222 -6662 132306 -6426
rect 132542 -6662 132574 -6426
rect 131954 -7654 132574 -6662
rect 151954 -7066 152574 33058
rect 160510 4045 160570 319363
rect 160794 282454 161414 321898
rect 160794 282218 160826 282454
rect 161382 282218 161414 282454
rect 160794 282134 161414 282218
rect 160794 281898 160826 282134
rect 161382 281898 161414 282134
rect 160794 242454 161414 281898
rect 160794 242218 160826 242454
rect 161382 242218 161414 242454
rect 160794 242134 161414 242218
rect 160794 241898 160826 242134
rect 161382 241898 161414 242134
rect 160794 202454 161414 241898
rect 160794 202218 160826 202454
rect 161382 202218 161414 202454
rect 160794 202134 161414 202218
rect 160794 201898 160826 202134
rect 161382 201898 161414 202134
rect 160794 162454 161414 201898
rect 160794 162218 160826 162454
rect 161382 162218 161414 162454
rect 160794 162134 161414 162218
rect 160794 161898 160826 162134
rect 161382 161898 161414 162134
rect 160794 122454 161414 161898
rect 160794 122218 160826 122454
rect 161062 122218 161146 122454
rect 161382 122218 161414 122454
rect 160794 122134 161414 122218
rect 160794 121898 160826 122134
rect 161062 121898 161146 122134
rect 161382 121898 161414 122134
rect 160794 82454 161414 121898
rect 160794 82218 160826 82454
rect 161062 82218 161146 82454
rect 161382 82218 161414 82454
rect 160794 82134 161414 82218
rect 160794 81898 160826 82134
rect 161062 81898 161146 82134
rect 161382 81898 161414 82134
rect 160794 42454 161414 81898
rect 160794 42218 160826 42454
rect 161062 42218 161146 42454
rect 161382 42218 161414 42454
rect 160794 42134 161414 42218
rect 160794 41898 160826 42134
rect 161062 41898 161146 42134
rect 161382 41898 161414 42134
rect 160507 4044 160573 4045
rect 160507 3980 160508 4044
rect 160572 3980 160573 4044
rect 160507 3979 160573 3980
rect 160794 2454 161414 41898
rect 160794 2218 160826 2454
rect 161062 2218 161146 2454
rect 161382 2218 161414 2454
rect 160794 2134 161414 2218
rect 160794 1898 160826 2134
rect 161062 1898 161146 2134
rect 161382 1898 161414 2134
rect 160794 -346 161414 1898
rect 160794 -582 160826 -346
rect 161062 -582 161146 -346
rect 161382 -582 161414 -346
rect 160794 -666 161414 -582
rect 160794 -902 160826 -666
rect 161062 -902 161146 -666
rect 161382 -902 161414 -666
rect 160794 -1894 161414 -902
rect 164514 686174 165134 706202
rect 164514 685938 164546 686174
rect 164782 685938 164866 686174
rect 165102 685938 165134 686174
rect 164514 685854 165134 685938
rect 164514 685618 164546 685854
rect 164782 685618 164866 685854
rect 165102 685618 165134 685854
rect 164514 646174 165134 685618
rect 164514 645938 164546 646174
rect 164782 645938 164866 646174
rect 165102 645938 165134 646174
rect 164514 645854 165134 645938
rect 164514 645618 164546 645854
rect 164782 645618 164866 645854
rect 165102 645618 165134 645854
rect 164514 606174 165134 645618
rect 164514 605938 164546 606174
rect 164782 605938 164866 606174
rect 165102 605938 165134 606174
rect 164514 605854 165134 605938
rect 164514 605618 164546 605854
rect 164782 605618 164866 605854
rect 165102 605618 165134 605854
rect 164514 566174 165134 605618
rect 164514 565938 164546 566174
rect 164782 565938 164866 566174
rect 165102 565938 165134 566174
rect 164514 565854 165134 565938
rect 164514 565618 164546 565854
rect 164782 565618 164866 565854
rect 165102 565618 165134 565854
rect 164514 526174 165134 565618
rect 164514 525938 164546 526174
rect 164782 525938 164866 526174
rect 165102 525938 165134 526174
rect 164514 525854 165134 525938
rect 164514 525618 164546 525854
rect 164782 525618 164866 525854
rect 165102 525618 165134 525854
rect 164514 486174 165134 525618
rect 164514 485938 164546 486174
rect 164782 485938 164866 486174
rect 165102 485938 165134 486174
rect 164514 485854 165134 485938
rect 164514 485618 164546 485854
rect 164782 485618 164866 485854
rect 165102 485618 165134 485854
rect 164514 446174 165134 485618
rect 164514 445938 164546 446174
rect 164782 445938 164866 446174
rect 165102 445938 165134 446174
rect 164514 445854 165134 445938
rect 164514 445618 164546 445854
rect 164782 445618 164866 445854
rect 165102 445618 165134 445854
rect 164514 406174 165134 445618
rect 164514 405938 164546 406174
rect 164782 405938 164866 406174
rect 165102 405938 165134 406174
rect 164514 405854 165134 405938
rect 164514 405618 164546 405854
rect 164782 405618 164866 405854
rect 165102 405618 165134 405854
rect 164514 366174 165134 405618
rect 164514 365938 164546 366174
rect 164782 365938 164866 366174
rect 165102 365938 165134 366174
rect 164514 365854 165134 365938
rect 164514 365618 164546 365854
rect 164782 365618 164866 365854
rect 165102 365618 165134 365854
rect 164514 326174 165134 365618
rect 164514 325938 164546 326174
rect 164782 325938 164866 326174
rect 165102 325938 165134 326174
rect 164514 325854 165134 325938
rect 164514 325618 164546 325854
rect 164782 325618 164866 325854
rect 165102 325618 165134 325854
rect 164514 286174 165134 325618
rect 164514 285938 164546 286174
rect 164782 285938 164866 286174
rect 165102 285938 165134 286174
rect 164514 285854 165134 285938
rect 164514 285618 164546 285854
rect 164782 285618 164866 285854
rect 165102 285618 165134 285854
rect 164514 246174 165134 285618
rect 164514 245938 164546 246174
rect 164782 245938 164866 246174
rect 165102 245938 165134 246174
rect 164514 245854 165134 245938
rect 164514 245618 164546 245854
rect 164782 245618 164866 245854
rect 165102 245618 165134 245854
rect 164514 206174 165134 245618
rect 164514 205938 164546 206174
rect 164782 205938 164866 206174
rect 165102 205938 165134 206174
rect 164514 205854 165134 205938
rect 164514 205618 164546 205854
rect 164782 205618 164866 205854
rect 165102 205618 165134 205854
rect 164514 166174 165134 205618
rect 164514 165938 164546 166174
rect 164782 165938 164866 166174
rect 165102 165938 165134 166174
rect 164514 165854 165134 165938
rect 164514 165618 164546 165854
rect 164782 165618 164866 165854
rect 165102 165618 165134 165854
rect 164514 126174 165134 165618
rect 164514 125938 164546 126174
rect 164782 125938 164866 126174
rect 165102 125938 165134 126174
rect 164514 125854 165134 125938
rect 164514 125618 164546 125854
rect 164782 125618 164866 125854
rect 165102 125618 165134 125854
rect 164514 86174 165134 125618
rect 164514 85938 164546 86174
rect 164782 85938 164866 86174
rect 165102 85938 165134 86174
rect 164514 85854 165134 85938
rect 164514 85618 164546 85854
rect 164782 85618 164866 85854
rect 165102 85618 165134 85854
rect 164514 46174 165134 85618
rect 164514 45938 164546 46174
rect 164782 45938 164866 46174
rect 165102 45938 165134 46174
rect 164514 45854 165134 45938
rect 164514 45618 164546 45854
rect 164782 45618 164866 45854
rect 165102 45618 165134 45854
rect 164514 6174 165134 45618
rect 164514 5938 164546 6174
rect 164782 5938 164866 6174
rect 165102 5938 165134 6174
rect 164514 5854 165134 5938
rect 164514 5618 164546 5854
rect 164782 5618 164866 5854
rect 165102 5618 165134 5854
rect 164514 -2266 165134 5618
rect 164514 -2502 164546 -2266
rect 164782 -2502 164866 -2266
rect 165102 -2502 165134 -2266
rect 164514 -2586 165134 -2502
rect 164514 -2822 164546 -2586
rect 164782 -2822 164866 -2586
rect 165102 -2822 165134 -2586
rect 164514 -3814 165134 -2822
rect 168234 689894 168854 708122
rect 168234 689658 168266 689894
rect 168502 689658 168586 689894
rect 168822 689658 168854 689894
rect 168234 689574 168854 689658
rect 168234 689338 168266 689574
rect 168502 689338 168586 689574
rect 168822 689338 168854 689574
rect 168234 649894 168854 689338
rect 168234 649658 168266 649894
rect 168502 649658 168586 649894
rect 168822 649658 168854 649894
rect 168234 649574 168854 649658
rect 168234 649338 168266 649574
rect 168502 649338 168586 649574
rect 168822 649338 168854 649574
rect 168234 609894 168854 649338
rect 168234 609658 168266 609894
rect 168502 609658 168586 609894
rect 168822 609658 168854 609894
rect 168234 609574 168854 609658
rect 168234 609338 168266 609574
rect 168502 609338 168586 609574
rect 168822 609338 168854 609574
rect 168234 569894 168854 609338
rect 168234 569658 168266 569894
rect 168502 569658 168586 569894
rect 168822 569658 168854 569894
rect 168234 569574 168854 569658
rect 168234 569338 168266 569574
rect 168502 569338 168586 569574
rect 168822 569338 168854 569574
rect 168234 529894 168854 569338
rect 168234 529658 168266 529894
rect 168502 529658 168586 529894
rect 168822 529658 168854 529894
rect 168234 529574 168854 529658
rect 168234 529338 168266 529574
rect 168502 529338 168586 529574
rect 168822 529338 168854 529574
rect 168234 489894 168854 529338
rect 168234 489658 168266 489894
rect 168502 489658 168586 489894
rect 168822 489658 168854 489894
rect 168234 489574 168854 489658
rect 168234 489338 168266 489574
rect 168502 489338 168586 489574
rect 168822 489338 168854 489574
rect 168234 449894 168854 489338
rect 168234 449658 168266 449894
rect 168502 449658 168586 449894
rect 168822 449658 168854 449894
rect 168234 449574 168854 449658
rect 168234 449338 168266 449574
rect 168502 449338 168586 449574
rect 168822 449338 168854 449574
rect 168234 409894 168854 449338
rect 168234 409658 168266 409894
rect 168502 409658 168586 409894
rect 168822 409658 168854 409894
rect 168234 409574 168854 409658
rect 168234 409338 168266 409574
rect 168502 409338 168586 409574
rect 168822 409338 168854 409574
rect 168234 369894 168854 409338
rect 168234 369658 168266 369894
rect 168502 369658 168586 369894
rect 168822 369658 168854 369894
rect 168234 369574 168854 369658
rect 168234 369338 168266 369574
rect 168502 369338 168586 369574
rect 168822 369338 168854 369574
rect 168234 329894 168854 369338
rect 168234 329658 168266 329894
rect 168502 329658 168586 329894
rect 168822 329658 168854 329894
rect 168234 329574 168854 329658
rect 168234 329338 168266 329574
rect 168502 329338 168586 329574
rect 168822 329338 168854 329574
rect 168234 289894 168854 329338
rect 171954 693614 172574 710042
rect 191954 711558 192574 711590
rect 191954 711322 191986 711558
rect 192222 711322 192306 711558
rect 192542 711322 192574 711558
rect 191954 711238 192574 711322
rect 191954 711002 191986 711238
rect 192222 711002 192306 711238
rect 192542 711002 192574 711238
rect 188234 709638 188854 709670
rect 188234 709402 188266 709638
rect 188502 709402 188586 709638
rect 188822 709402 188854 709638
rect 188234 709318 188854 709402
rect 188234 709082 188266 709318
rect 188502 709082 188586 709318
rect 188822 709082 188854 709318
rect 184514 707718 185134 707750
rect 184514 707482 184546 707718
rect 184782 707482 184866 707718
rect 185102 707482 185134 707718
rect 184514 707398 185134 707482
rect 184514 707162 184546 707398
rect 184782 707162 184866 707398
rect 185102 707162 185134 707398
rect 171954 693378 171986 693614
rect 172222 693378 172306 693614
rect 172542 693378 172574 693614
rect 171954 693294 172574 693378
rect 171954 693058 171986 693294
rect 172222 693058 172306 693294
rect 172542 693058 172574 693294
rect 171954 653614 172574 693058
rect 171954 653378 171986 653614
rect 172222 653378 172306 653614
rect 172542 653378 172574 653614
rect 171954 653294 172574 653378
rect 171954 653058 171986 653294
rect 172222 653058 172306 653294
rect 172542 653058 172574 653294
rect 171954 613614 172574 653058
rect 171954 613378 171986 613614
rect 172222 613378 172306 613614
rect 172542 613378 172574 613614
rect 171954 613294 172574 613378
rect 171954 613058 171986 613294
rect 172222 613058 172306 613294
rect 172542 613058 172574 613294
rect 171954 573614 172574 613058
rect 171954 573378 171986 573614
rect 172222 573378 172306 573614
rect 172542 573378 172574 573614
rect 171954 573294 172574 573378
rect 171954 573058 171986 573294
rect 172222 573058 172306 573294
rect 172542 573058 172574 573294
rect 171954 533614 172574 573058
rect 171954 533378 171986 533614
rect 172222 533378 172306 533614
rect 172542 533378 172574 533614
rect 171954 533294 172574 533378
rect 171954 533058 171986 533294
rect 172222 533058 172306 533294
rect 172542 533058 172574 533294
rect 171954 493614 172574 533058
rect 171954 493378 171986 493614
rect 172222 493378 172306 493614
rect 172542 493378 172574 493614
rect 171954 493294 172574 493378
rect 171954 493058 171986 493294
rect 172222 493058 172306 493294
rect 172542 493058 172574 493294
rect 171954 453614 172574 493058
rect 171954 453378 171986 453614
rect 172222 453378 172306 453614
rect 172542 453378 172574 453614
rect 171954 453294 172574 453378
rect 171954 453058 171986 453294
rect 172222 453058 172306 453294
rect 172542 453058 172574 453294
rect 171954 413614 172574 453058
rect 171954 413378 171986 413614
rect 172222 413378 172306 413614
rect 172542 413378 172574 413614
rect 171954 413294 172574 413378
rect 171954 413058 171986 413294
rect 172222 413058 172306 413294
rect 172542 413058 172574 413294
rect 171954 373614 172574 413058
rect 171954 373378 171986 373614
rect 172222 373378 172306 373614
rect 172542 373378 172574 373614
rect 171954 373294 172574 373378
rect 171954 373058 171986 373294
rect 172222 373058 172306 373294
rect 172542 373058 172574 373294
rect 171954 333614 172574 373058
rect 171954 333378 171986 333614
rect 172222 333378 172306 333614
rect 172542 333378 172574 333614
rect 171954 333294 172574 333378
rect 171954 333058 171986 333294
rect 172222 333058 172306 333294
rect 172542 333058 172574 333294
rect 169707 319428 169773 319429
rect 169707 319364 169708 319428
rect 169772 319364 169773 319428
rect 169707 319363 169773 319364
rect 168234 289658 168266 289894
rect 168502 289658 168586 289894
rect 168822 289658 168854 289894
rect 168234 289574 168854 289658
rect 168234 289338 168266 289574
rect 168502 289338 168586 289574
rect 168822 289338 168854 289574
rect 168234 249894 168854 289338
rect 168234 249658 168266 249894
rect 168502 249658 168586 249894
rect 168822 249658 168854 249894
rect 168234 249574 168854 249658
rect 168234 249338 168266 249574
rect 168502 249338 168586 249574
rect 168822 249338 168854 249574
rect 168234 209894 168854 249338
rect 168234 209658 168266 209894
rect 168502 209658 168586 209894
rect 168822 209658 168854 209894
rect 168234 209574 168854 209658
rect 168234 209338 168266 209574
rect 168502 209338 168586 209574
rect 168822 209338 168854 209574
rect 168234 169894 168854 209338
rect 168234 169658 168266 169894
rect 168502 169658 168586 169894
rect 168822 169658 168854 169894
rect 168234 169574 168854 169658
rect 168234 169338 168266 169574
rect 168502 169338 168586 169574
rect 168822 169338 168854 169574
rect 168234 129894 168854 169338
rect 168234 129658 168266 129894
rect 168502 129658 168586 129894
rect 168822 129658 168854 129894
rect 168234 129574 168854 129658
rect 168234 129338 168266 129574
rect 168502 129338 168586 129574
rect 168822 129338 168854 129574
rect 168234 89894 168854 129338
rect 168234 89658 168266 89894
rect 168502 89658 168586 89894
rect 168822 89658 168854 89894
rect 168234 89574 168854 89658
rect 168234 89338 168266 89574
rect 168502 89338 168586 89574
rect 168822 89338 168854 89574
rect 168234 49894 168854 89338
rect 168234 49658 168266 49894
rect 168502 49658 168586 49894
rect 168822 49658 168854 49894
rect 168234 49574 168854 49658
rect 168234 49338 168266 49574
rect 168502 49338 168586 49574
rect 168822 49338 168854 49574
rect 168234 9894 168854 49338
rect 168234 9658 168266 9894
rect 168502 9658 168586 9894
rect 168822 9658 168854 9894
rect 168234 9574 168854 9658
rect 168234 9338 168266 9574
rect 168502 9338 168586 9574
rect 168822 9338 168854 9574
rect 168234 -4186 168854 9338
rect 169710 3773 169770 319363
rect 171954 293614 172574 333058
rect 180794 705798 181414 705830
rect 180794 705562 180826 705798
rect 181062 705562 181146 705798
rect 181382 705562 181414 705798
rect 180794 705478 181414 705562
rect 180794 705242 180826 705478
rect 181062 705242 181146 705478
rect 181382 705242 181414 705478
rect 180794 662454 181414 705242
rect 180794 662218 180826 662454
rect 181062 662218 181146 662454
rect 181382 662218 181414 662454
rect 180794 662134 181414 662218
rect 180794 661898 180826 662134
rect 181062 661898 181146 662134
rect 181382 661898 181414 662134
rect 180794 622454 181414 661898
rect 180794 622218 180826 622454
rect 181062 622218 181146 622454
rect 181382 622218 181414 622454
rect 180794 622134 181414 622218
rect 180794 621898 180826 622134
rect 181062 621898 181146 622134
rect 181382 621898 181414 622134
rect 180794 582454 181414 621898
rect 180794 582218 180826 582454
rect 181062 582218 181146 582454
rect 181382 582218 181414 582454
rect 180794 582134 181414 582218
rect 180794 581898 180826 582134
rect 181062 581898 181146 582134
rect 181382 581898 181414 582134
rect 180794 542454 181414 581898
rect 180794 542218 180826 542454
rect 181062 542218 181146 542454
rect 181382 542218 181414 542454
rect 180794 542134 181414 542218
rect 180794 541898 180826 542134
rect 181062 541898 181146 542134
rect 181382 541898 181414 542134
rect 180794 502454 181414 541898
rect 180794 502218 180826 502454
rect 181062 502218 181146 502454
rect 181382 502218 181414 502454
rect 180794 502134 181414 502218
rect 180794 501898 180826 502134
rect 181062 501898 181146 502134
rect 181382 501898 181414 502134
rect 180794 462454 181414 501898
rect 180794 462218 180826 462454
rect 181062 462218 181146 462454
rect 181382 462218 181414 462454
rect 180794 462134 181414 462218
rect 180794 461898 180826 462134
rect 181062 461898 181146 462134
rect 181382 461898 181414 462134
rect 180794 422454 181414 461898
rect 180794 422218 180826 422454
rect 181062 422218 181146 422454
rect 181382 422218 181414 422454
rect 180794 422134 181414 422218
rect 180794 421898 180826 422134
rect 181062 421898 181146 422134
rect 181382 421898 181414 422134
rect 180794 382454 181414 421898
rect 180794 382218 180826 382454
rect 181062 382218 181146 382454
rect 181382 382218 181414 382454
rect 180794 382134 181414 382218
rect 180794 381898 180826 382134
rect 181062 381898 181146 382134
rect 181382 381898 181414 382134
rect 180794 342454 181414 381898
rect 180794 342218 180826 342454
rect 181062 342218 181146 342454
rect 181382 342218 181414 342454
rect 180794 342134 181414 342218
rect 180794 341898 180826 342134
rect 181062 341898 181146 342134
rect 181382 341898 181414 342134
rect 179459 319428 179525 319429
rect 179459 319364 179460 319428
rect 179524 319364 179525 319428
rect 179459 319363 179525 319364
rect 171954 293378 171986 293614
rect 172222 293378 172306 293614
rect 172542 293378 172574 293614
rect 171954 293294 172574 293378
rect 171954 293058 171986 293294
rect 172222 293058 172306 293294
rect 172542 293058 172574 293294
rect 171954 253614 172574 293058
rect 171954 253378 171986 253614
rect 172222 253378 172306 253614
rect 172542 253378 172574 253614
rect 171954 253294 172574 253378
rect 171954 253058 171986 253294
rect 172222 253058 172306 253294
rect 172542 253058 172574 253294
rect 171954 213614 172574 253058
rect 171954 213378 171986 213614
rect 172222 213378 172306 213614
rect 172542 213378 172574 213614
rect 171954 213294 172574 213378
rect 171954 213058 171986 213294
rect 172222 213058 172306 213294
rect 172542 213058 172574 213294
rect 171954 173614 172574 213058
rect 171954 173378 171986 173614
rect 172222 173378 172306 173614
rect 172542 173378 172574 173614
rect 171954 173294 172574 173378
rect 171954 173058 171986 173294
rect 172222 173058 172306 173294
rect 172542 173058 172574 173294
rect 171954 133614 172574 173058
rect 171954 133378 171986 133614
rect 172222 133378 172306 133614
rect 172542 133378 172574 133614
rect 171954 133294 172574 133378
rect 171954 133058 171986 133294
rect 172222 133058 172306 133294
rect 172542 133058 172574 133294
rect 171954 93614 172574 133058
rect 171954 93378 171986 93614
rect 172222 93378 172306 93614
rect 172542 93378 172574 93614
rect 171954 93294 172574 93378
rect 171954 93058 171986 93294
rect 172222 93058 172306 93294
rect 172542 93058 172574 93294
rect 171954 53614 172574 93058
rect 171954 53378 171986 53614
rect 172222 53378 172306 53614
rect 172542 53378 172574 53614
rect 171954 53294 172574 53378
rect 171954 53058 171986 53294
rect 172222 53058 172306 53294
rect 172542 53058 172574 53294
rect 171954 13614 172574 53058
rect 171954 13378 171986 13614
rect 172222 13378 172306 13614
rect 172542 13378 172574 13614
rect 171954 13294 172574 13378
rect 171954 13058 171986 13294
rect 172222 13058 172306 13294
rect 172542 13058 172574 13294
rect 169707 3772 169773 3773
rect 169707 3708 169708 3772
rect 169772 3708 169773 3772
rect 169707 3707 169773 3708
rect 168234 -4422 168266 -4186
rect 168502 -4422 168586 -4186
rect 168822 -4422 168854 -4186
rect 168234 -4506 168854 -4422
rect 168234 -4742 168266 -4506
rect 168502 -4742 168586 -4506
rect 168822 -4742 168854 -4506
rect 168234 -5734 168854 -4742
rect 151954 -7302 151986 -7066
rect 152222 -7302 152306 -7066
rect 152542 -7302 152574 -7066
rect 151954 -7386 152574 -7302
rect 151954 -7622 151986 -7386
rect 152222 -7622 152306 -7386
rect 152542 -7622 152574 -7386
rect 151954 -7654 152574 -7622
rect 171954 -6106 172574 13058
rect 179462 3909 179522 319363
rect 180794 302454 181414 341898
rect 180794 302218 180826 302454
rect 181382 302218 181414 302454
rect 180794 302134 181414 302218
rect 180794 301898 180826 302134
rect 181382 301898 181414 302134
rect 180794 262454 181414 301898
rect 180794 262218 180826 262454
rect 181382 262218 181414 262454
rect 180794 262134 181414 262218
rect 180794 261898 180826 262134
rect 181382 261898 181414 262134
rect 180794 222454 181414 261898
rect 180794 222218 180826 222454
rect 181382 222218 181414 222454
rect 180794 222134 181414 222218
rect 180794 221898 180826 222134
rect 181382 221898 181414 222134
rect 180794 182454 181414 221898
rect 180794 182218 180826 182454
rect 181382 182218 181414 182454
rect 180794 182134 181414 182218
rect 180794 181898 180826 182134
rect 181382 181898 181414 182134
rect 180794 142454 181414 181898
rect 180794 142218 180826 142454
rect 181382 142218 181414 142454
rect 180794 142134 181414 142218
rect 180794 141898 180826 142134
rect 181382 141898 181414 142134
rect 180794 102454 181414 141898
rect 180794 102218 180826 102454
rect 181062 102218 181146 102454
rect 181382 102218 181414 102454
rect 180794 102134 181414 102218
rect 180794 101898 180826 102134
rect 181062 101898 181146 102134
rect 181382 101898 181414 102134
rect 180794 62454 181414 101898
rect 180794 62218 180826 62454
rect 181062 62218 181146 62454
rect 181382 62218 181414 62454
rect 180794 62134 181414 62218
rect 180794 61898 180826 62134
rect 181062 61898 181146 62134
rect 181382 61898 181414 62134
rect 180794 22454 181414 61898
rect 180794 22218 180826 22454
rect 181062 22218 181146 22454
rect 181382 22218 181414 22454
rect 180794 22134 181414 22218
rect 180794 21898 180826 22134
rect 181062 21898 181146 22134
rect 181382 21898 181414 22134
rect 179459 3908 179525 3909
rect 179459 3844 179460 3908
rect 179524 3844 179525 3908
rect 179459 3843 179525 3844
rect 180794 -1306 181414 21898
rect 180794 -1542 180826 -1306
rect 181062 -1542 181146 -1306
rect 181382 -1542 181414 -1306
rect 180794 -1626 181414 -1542
rect 180794 -1862 180826 -1626
rect 181062 -1862 181146 -1626
rect 181382 -1862 181414 -1626
rect 180794 -1894 181414 -1862
rect 184514 666174 185134 707162
rect 184514 665938 184546 666174
rect 184782 665938 184866 666174
rect 185102 665938 185134 666174
rect 184514 665854 185134 665938
rect 184514 665618 184546 665854
rect 184782 665618 184866 665854
rect 185102 665618 185134 665854
rect 184514 626174 185134 665618
rect 184514 625938 184546 626174
rect 184782 625938 184866 626174
rect 185102 625938 185134 626174
rect 184514 625854 185134 625938
rect 184514 625618 184546 625854
rect 184782 625618 184866 625854
rect 185102 625618 185134 625854
rect 184514 586174 185134 625618
rect 184514 585938 184546 586174
rect 184782 585938 184866 586174
rect 185102 585938 185134 586174
rect 184514 585854 185134 585938
rect 184514 585618 184546 585854
rect 184782 585618 184866 585854
rect 185102 585618 185134 585854
rect 184514 546174 185134 585618
rect 184514 545938 184546 546174
rect 184782 545938 184866 546174
rect 185102 545938 185134 546174
rect 184514 545854 185134 545938
rect 184514 545618 184546 545854
rect 184782 545618 184866 545854
rect 185102 545618 185134 545854
rect 184514 506174 185134 545618
rect 184514 505938 184546 506174
rect 184782 505938 184866 506174
rect 185102 505938 185134 506174
rect 184514 505854 185134 505938
rect 184514 505618 184546 505854
rect 184782 505618 184866 505854
rect 185102 505618 185134 505854
rect 184514 466174 185134 505618
rect 184514 465938 184546 466174
rect 184782 465938 184866 466174
rect 185102 465938 185134 466174
rect 184514 465854 185134 465938
rect 184514 465618 184546 465854
rect 184782 465618 184866 465854
rect 185102 465618 185134 465854
rect 184514 426174 185134 465618
rect 184514 425938 184546 426174
rect 184782 425938 184866 426174
rect 185102 425938 185134 426174
rect 184514 425854 185134 425938
rect 184514 425618 184546 425854
rect 184782 425618 184866 425854
rect 185102 425618 185134 425854
rect 184514 386174 185134 425618
rect 184514 385938 184546 386174
rect 184782 385938 184866 386174
rect 185102 385938 185134 386174
rect 184514 385854 185134 385938
rect 184514 385618 184546 385854
rect 184782 385618 184866 385854
rect 185102 385618 185134 385854
rect 184514 346174 185134 385618
rect 184514 345938 184546 346174
rect 184782 345938 184866 346174
rect 185102 345938 185134 346174
rect 184514 345854 185134 345938
rect 184514 345618 184546 345854
rect 184782 345618 184866 345854
rect 185102 345618 185134 345854
rect 184514 306174 185134 345618
rect 184514 305938 184546 306174
rect 184782 305938 184866 306174
rect 185102 305938 185134 306174
rect 184514 305854 185134 305938
rect 184514 305618 184546 305854
rect 184782 305618 184866 305854
rect 185102 305618 185134 305854
rect 184514 266174 185134 305618
rect 184514 265938 184546 266174
rect 184782 265938 184866 266174
rect 185102 265938 185134 266174
rect 184514 265854 185134 265938
rect 184514 265618 184546 265854
rect 184782 265618 184866 265854
rect 185102 265618 185134 265854
rect 184514 226174 185134 265618
rect 184514 225938 184546 226174
rect 184782 225938 184866 226174
rect 185102 225938 185134 226174
rect 184514 225854 185134 225938
rect 184514 225618 184546 225854
rect 184782 225618 184866 225854
rect 185102 225618 185134 225854
rect 184514 186174 185134 225618
rect 184514 185938 184546 186174
rect 184782 185938 184866 186174
rect 185102 185938 185134 186174
rect 184514 185854 185134 185938
rect 184514 185618 184546 185854
rect 184782 185618 184866 185854
rect 185102 185618 185134 185854
rect 184514 146174 185134 185618
rect 184514 145938 184546 146174
rect 184782 145938 184866 146174
rect 185102 145938 185134 146174
rect 184514 145854 185134 145938
rect 184514 145618 184546 145854
rect 184782 145618 184866 145854
rect 185102 145618 185134 145854
rect 184514 106174 185134 145618
rect 184514 105938 184546 106174
rect 184782 105938 184866 106174
rect 185102 105938 185134 106174
rect 184514 105854 185134 105938
rect 184514 105618 184546 105854
rect 184782 105618 184866 105854
rect 185102 105618 185134 105854
rect 184514 66174 185134 105618
rect 184514 65938 184546 66174
rect 184782 65938 184866 66174
rect 185102 65938 185134 66174
rect 184514 65854 185134 65938
rect 184514 65618 184546 65854
rect 184782 65618 184866 65854
rect 185102 65618 185134 65854
rect 184514 26174 185134 65618
rect 184514 25938 184546 26174
rect 184782 25938 184866 26174
rect 185102 25938 185134 26174
rect 184514 25854 185134 25938
rect 184514 25618 184546 25854
rect 184782 25618 184866 25854
rect 185102 25618 185134 25854
rect 184514 -3226 185134 25618
rect 184514 -3462 184546 -3226
rect 184782 -3462 184866 -3226
rect 185102 -3462 185134 -3226
rect 184514 -3546 185134 -3462
rect 184514 -3782 184546 -3546
rect 184782 -3782 184866 -3546
rect 185102 -3782 185134 -3546
rect 184514 -3814 185134 -3782
rect 188234 669894 188854 709082
rect 188234 669658 188266 669894
rect 188502 669658 188586 669894
rect 188822 669658 188854 669894
rect 188234 669574 188854 669658
rect 188234 669338 188266 669574
rect 188502 669338 188586 669574
rect 188822 669338 188854 669574
rect 188234 629894 188854 669338
rect 188234 629658 188266 629894
rect 188502 629658 188586 629894
rect 188822 629658 188854 629894
rect 188234 629574 188854 629658
rect 188234 629338 188266 629574
rect 188502 629338 188586 629574
rect 188822 629338 188854 629574
rect 188234 589894 188854 629338
rect 188234 589658 188266 589894
rect 188502 589658 188586 589894
rect 188822 589658 188854 589894
rect 188234 589574 188854 589658
rect 188234 589338 188266 589574
rect 188502 589338 188586 589574
rect 188822 589338 188854 589574
rect 188234 549894 188854 589338
rect 188234 549658 188266 549894
rect 188502 549658 188586 549894
rect 188822 549658 188854 549894
rect 188234 549574 188854 549658
rect 188234 549338 188266 549574
rect 188502 549338 188586 549574
rect 188822 549338 188854 549574
rect 188234 509894 188854 549338
rect 188234 509658 188266 509894
rect 188502 509658 188586 509894
rect 188822 509658 188854 509894
rect 188234 509574 188854 509658
rect 188234 509338 188266 509574
rect 188502 509338 188586 509574
rect 188822 509338 188854 509574
rect 188234 469894 188854 509338
rect 188234 469658 188266 469894
rect 188502 469658 188586 469894
rect 188822 469658 188854 469894
rect 188234 469574 188854 469658
rect 188234 469338 188266 469574
rect 188502 469338 188586 469574
rect 188822 469338 188854 469574
rect 188234 429894 188854 469338
rect 188234 429658 188266 429894
rect 188502 429658 188586 429894
rect 188822 429658 188854 429894
rect 188234 429574 188854 429658
rect 188234 429338 188266 429574
rect 188502 429338 188586 429574
rect 188822 429338 188854 429574
rect 188234 389894 188854 429338
rect 188234 389658 188266 389894
rect 188502 389658 188586 389894
rect 188822 389658 188854 389894
rect 188234 389574 188854 389658
rect 188234 389338 188266 389574
rect 188502 389338 188586 389574
rect 188822 389338 188854 389574
rect 188234 349894 188854 389338
rect 188234 349658 188266 349894
rect 188502 349658 188586 349894
rect 188822 349658 188854 349894
rect 188234 349574 188854 349658
rect 188234 349338 188266 349574
rect 188502 349338 188586 349574
rect 188822 349338 188854 349574
rect 188234 309894 188854 349338
rect 188234 309658 188266 309894
rect 188502 309658 188586 309894
rect 188822 309658 188854 309894
rect 188234 309574 188854 309658
rect 188234 309338 188266 309574
rect 188502 309338 188586 309574
rect 188822 309338 188854 309574
rect 188234 269894 188854 309338
rect 188234 269658 188266 269894
rect 188502 269658 188586 269894
rect 188822 269658 188854 269894
rect 188234 269574 188854 269658
rect 188234 269338 188266 269574
rect 188502 269338 188586 269574
rect 188822 269338 188854 269574
rect 188234 229894 188854 269338
rect 188234 229658 188266 229894
rect 188502 229658 188586 229894
rect 188822 229658 188854 229894
rect 188234 229574 188854 229658
rect 188234 229338 188266 229574
rect 188502 229338 188586 229574
rect 188822 229338 188854 229574
rect 188234 189894 188854 229338
rect 188234 189658 188266 189894
rect 188502 189658 188586 189894
rect 188822 189658 188854 189894
rect 188234 189574 188854 189658
rect 188234 189338 188266 189574
rect 188502 189338 188586 189574
rect 188822 189338 188854 189574
rect 188234 149894 188854 189338
rect 188234 149658 188266 149894
rect 188502 149658 188586 149894
rect 188822 149658 188854 149894
rect 188234 149574 188854 149658
rect 188234 149338 188266 149574
rect 188502 149338 188586 149574
rect 188822 149338 188854 149574
rect 188234 109894 188854 149338
rect 188234 109658 188266 109894
rect 188502 109658 188586 109894
rect 188822 109658 188854 109894
rect 188234 109574 188854 109658
rect 188234 109338 188266 109574
rect 188502 109338 188586 109574
rect 188822 109338 188854 109574
rect 188234 69894 188854 109338
rect 188234 69658 188266 69894
rect 188502 69658 188586 69894
rect 188822 69658 188854 69894
rect 188234 69574 188854 69658
rect 188234 69338 188266 69574
rect 188502 69338 188586 69574
rect 188822 69338 188854 69574
rect 188234 29894 188854 69338
rect 188234 29658 188266 29894
rect 188502 29658 188586 29894
rect 188822 29658 188854 29894
rect 188234 29574 188854 29658
rect 188234 29338 188266 29574
rect 188502 29338 188586 29574
rect 188822 29338 188854 29574
rect 188234 -5146 188854 29338
rect 188234 -5382 188266 -5146
rect 188502 -5382 188586 -5146
rect 188822 -5382 188854 -5146
rect 188234 -5466 188854 -5382
rect 188234 -5702 188266 -5466
rect 188502 -5702 188586 -5466
rect 188822 -5702 188854 -5466
rect 188234 -5734 188854 -5702
rect 191954 673614 192574 711002
rect 211954 710598 212574 711590
rect 211954 710362 211986 710598
rect 212222 710362 212306 710598
rect 212542 710362 212574 710598
rect 211954 710278 212574 710362
rect 211954 710042 211986 710278
rect 212222 710042 212306 710278
rect 212542 710042 212574 710278
rect 208234 708678 208854 709670
rect 208234 708442 208266 708678
rect 208502 708442 208586 708678
rect 208822 708442 208854 708678
rect 208234 708358 208854 708442
rect 208234 708122 208266 708358
rect 208502 708122 208586 708358
rect 208822 708122 208854 708358
rect 204514 706758 205134 707750
rect 204514 706522 204546 706758
rect 204782 706522 204866 706758
rect 205102 706522 205134 706758
rect 204514 706438 205134 706522
rect 204514 706202 204546 706438
rect 204782 706202 204866 706438
rect 205102 706202 205134 706438
rect 191954 673378 191986 673614
rect 192222 673378 192306 673614
rect 192542 673378 192574 673614
rect 191954 673294 192574 673378
rect 191954 673058 191986 673294
rect 192222 673058 192306 673294
rect 192542 673058 192574 673294
rect 191954 633614 192574 673058
rect 191954 633378 191986 633614
rect 192222 633378 192306 633614
rect 192542 633378 192574 633614
rect 191954 633294 192574 633378
rect 191954 633058 191986 633294
rect 192222 633058 192306 633294
rect 192542 633058 192574 633294
rect 191954 593614 192574 633058
rect 191954 593378 191986 593614
rect 192222 593378 192306 593614
rect 192542 593378 192574 593614
rect 191954 593294 192574 593378
rect 191954 593058 191986 593294
rect 192222 593058 192306 593294
rect 192542 593058 192574 593294
rect 191954 553614 192574 593058
rect 191954 553378 191986 553614
rect 192222 553378 192306 553614
rect 192542 553378 192574 553614
rect 191954 553294 192574 553378
rect 191954 553058 191986 553294
rect 192222 553058 192306 553294
rect 192542 553058 192574 553294
rect 191954 513614 192574 553058
rect 191954 513378 191986 513614
rect 192222 513378 192306 513614
rect 192542 513378 192574 513614
rect 191954 513294 192574 513378
rect 191954 513058 191986 513294
rect 192222 513058 192306 513294
rect 192542 513058 192574 513294
rect 191954 473614 192574 513058
rect 191954 473378 191986 473614
rect 192222 473378 192306 473614
rect 192542 473378 192574 473614
rect 191954 473294 192574 473378
rect 191954 473058 191986 473294
rect 192222 473058 192306 473294
rect 192542 473058 192574 473294
rect 191954 433614 192574 473058
rect 191954 433378 191986 433614
rect 192222 433378 192306 433614
rect 192542 433378 192574 433614
rect 191954 433294 192574 433378
rect 191954 433058 191986 433294
rect 192222 433058 192306 433294
rect 192542 433058 192574 433294
rect 191954 393614 192574 433058
rect 191954 393378 191986 393614
rect 192222 393378 192306 393614
rect 192542 393378 192574 393614
rect 191954 393294 192574 393378
rect 191954 393058 191986 393294
rect 192222 393058 192306 393294
rect 192542 393058 192574 393294
rect 191954 353614 192574 393058
rect 191954 353378 191986 353614
rect 192222 353378 192306 353614
rect 192542 353378 192574 353614
rect 191954 353294 192574 353378
rect 191954 353058 191986 353294
rect 192222 353058 192306 353294
rect 192542 353058 192574 353294
rect 191954 313614 192574 353058
rect 200794 704838 201414 705830
rect 200794 704602 200826 704838
rect 201062 704602 201146 704838
rect 201382 704602 201414 704838
rect 200794 704518 201414 704602
rect 200794 704282 200826 704518
rect 201062 704282 201146 704518
rect 201382 704282 201414 704518
rect 200794 682454 201414 704282
rect 200794 682218 200826 682454
rect 201062 682218 201146 682454
rect 201382 682218 201414 682454
rect 200794 682134 201414 682218
rect 200794 681898 200826 682134
rect 201062 681898 201146 682134
rect 201382 681898 201414 682134
rect 200794 642454 201414 681898
rect 200794 642218 200826 642454
rect 201062 642218 201146 642454
rect 201382 642218 201414 642454
rect 200794 642134 201414 642218
rect 200794 641898 200826 642134
rect 201062 641898 201146 642134
rect 201382 641898 201414 642134
rect 200794 602454 201414 641898
rect 200794 602218 200826 602454
rect 201062 602218 201146 602454
rect 201382 602218 201414 602454
rect 200794 602134 201414 602218
rect 200794 601898 200826 602134
rect 201062 601898 201146 602134
rect 201382 601898 201414 602134
rect 200794 562454 201414 601898
rect 200794 562218 200826 562454
rect 201062 562218 201146 562454
rect 201382 562218 201414 562454
rect 200794 562134 201414 562218
rect 200794 561898 200826 562134
rect 201062 561898 201146 562134
rect 201382 561898 201414 562134
rect 200794 522454 201414 561898
rect 200794 522218 200826 522454
rect 201062 522218 201146 522454
rect 201382 522218 201414 522454
rect 200794 522134 201414 522218
rect 200794 521898 200826 522134
rect 201062 521898 201146 522134
rect 201382 521898 201414 522134
rect 200794 482454 201414 521898
rect 200794 482218 200826 482454
rect 201062 482218 201146 482454
rect 201382 482218 201414 482454
rect 200794 482134 201414 482218
rect 200794 481898 200826 482134
rect 201062 481898 201146 482134
rect 201382 481898 201414 482134
rect 200794 442454 201414 481898
rect 200794 442218 200826 442454
rect 201062 442218 201146 442454
rect 201382 442218 201414 442454
rect 200794 442134 201414 442218
rect 200794 441898 200826 442134
rect 201062 441898 201146 442134
rect 201382 441898 201414 442134
rect 200794 402454 201414 441898
rect 200794 402218 200826 402454
rect 201062 402218 201146 402454
rect 201382 402218 201414 402454
rect 200794 402134 201414 402218
rect 200794 401898 200826 402134
rect 201062 401898 201146 402134
rect 201382 401898 201414 402134
rect 200794 362454 201414 401898
rect 200794 362218 200826 362454
rect 201062 362218 201146 362454
rect 201382 362218 201414 362454
rect 200794 362134 201414 362218
rect 200794 361898 200826 362134
rect 201062 361898 201146 362134
rect 201382 361898 201414 362134
rect 200794 322454 201414 361898
rect 200794 322218 200826 322454
rect 201062 322218 201146 322454
rect 201382 322218 201414 322454
rect 200794 322134 201414 322218
rect 200794 321898 200826 322134
rect 201062 321898 201146 322134
rect 201382 321898 201414 322134
rect 200251 319428 200317 319429
rect 200251 319364 200252 319428
rect 200316 319364 200317 319428
rect 200251 319363 200317 319364
rect 200254 319290 200314 319363
rect 191954 313378 191986 313614
rect 192222 313378 192306 313614
rect 192542 313378 192574 313614
rect 191954 313294 192574 313378
rect 191954 313058 191986 313294
rect 192222 313058 192306 313294
rect 192542 313058 192574 313294
rect 191954 273614 192574 313058
rect 191954 273378 191986 273614
rect 192222 273378 192306 273614
rect 192542 273378 192574 273614
rect 191954 273294 192574 273378
rect 191954 273058 191986 273294
rect 192222 273058 192306 273294
rect 192542 273058 192574 273294
rect 191954 233614 192574 273058
rect 191954 233378 191986 233614
rect 192222 233378 192306 233614
rect 192542 233378 192574 233614
rect 191954 233294 192574 233378
rect 191954 233058 191986 233294
rect 192222 233058 192306 233294
rect 192542 233058 192574 233294
rect 191954 193614 192574 233058
rect 191954 193378 191986 193614
rect 192222 193378 192306 193614
rect 192542 193378 192574 193614
rect 191954 193294 192574 193378
rect 191954 193058 191986 193294
rect 192222 193058 192306 193294
rect 192542 193058 192574 193294
rect 191954 153614 192574 193058
rect 191954 153378 191986 153614
rect 192222 153378 192306 153614
rect 192542 153378 192574 153614
rect 191954 153294 192574 153378
rect 191954 153058 191986 153294
rect 192222 153058 192306 153294
rect 192542 153058 192574 153294
rect 191954 113614 192574 153058
rect 191954 113378 191986 113614
rect 192222 113378 192306 113614
rect 192542 113378 192574 113614
rect 191954 113294 192574 113378
rect 191954 113058 191986 113294
rect 192222 113058 192306 113294
rect 192542 113058 192574 113294
rect 191954 73614 192574 113058
rect 191954 73378 191986 73614
rect 192222 73378 192306 73614
rect 192542 73378 192574 73614
rect 191954 73294 192574 73378
rect 191954 73058 191986 73294
rect 192222 73058 192306 73294
rect 192542 73058 192574 73294
rect 191954 33614 192574 73058
rect 191954 33378 191986 33614
rect 192222 33378 192306 33614
rect 192542 33378 192574 33614
rect 191954 33294 192574 33378
rect 191954 33058 191986 33294
rect 192222 33058 192306 33294
rect 192542 33058 192574 33294
rect 171954 -6342 171986 -6106
rect 172222 -6342 172306 -6106
rect 172542 -6342 172574 -6106
rect 171954 -6426 172574 -6342
rect 171954 -6662 171986 -6426
rect 172222 -6662 172306 -6426
rect 172542 -6662 172574 -6426
rect 171954 -7654 172574 -6662
rect 191954 -7066 192574 33058
rect 199886 319230 200314 319290
rect 199886 3637 199946 319230
rect 200794 282454 201414 321898
rect 200794 282218 200826 282454
rect 201382 282218 201414 282454
rect 200794 282134 201414 282218
rect 200794 281898 200826 282134
rect 201382 281898 201414 282134
rect 200794 242454 201414 281898
rect 200794 242218 200826 242454
rect 201382 242218 201414 242454
rect 200794 242134 201414 242218
rect 200794 241898 200826 242134
rect 201382 241898 201414 242134
rect 200794 202454 201414 241898
rect 200794 202218 200826 202454
rect 201382 202218 201414 202454
rect 200794 202134 201414 202218
rect 200794 201898 200826 202134
rect 201382 201898 201414 202134
rect 200794 162454 201414 201898
rect 200794 162218 200826 162454
rect 201382 162218 201414 162454
rect 200794 162134 201414 162218
rect 200794 161898 200826 162134
rect 201382 161898 201414 162134
rect 200794 122454 201414 161898
rect 200794 122218 200826 122454
rect 201062 122218 201146 122454
rect 201382 122218 201414 122454
rect 200794 122134 201414 122218
rect 200794 121898 200826 122134
rect 201062 121898 201146 122134
rect 201382 121898 201414 122134
rect 200794 82454 201414 121898
rect 200794 82218 200826 82454
rect 201062 82218 201146 82454
rect 201382 82218 201414 82454
rect 200794 82134 201414 82218
rect 200794 81898 200826 82134
rect 201062 81898 201146 82134
rect 201382 81898 201414 82134
rect 200794 42454 201414 81898
rect 200794 42218 200826 42454
rect 201062 42218 201146 42454
rect 201382 42218 201414 42454
rect 200794 42134 201414 42218
rect 200794 41898 200826 42134
rect 201062 41898 201146 42134
rect 201382 41898 201414 42134
rect 199883 3636 199949 3637
rect 199883 3572 199884 3636
rect 199948 3572 199949 3636
rect 199883 3571 199949 3572
rect 200794 2454 201414 41898
rect 200794 2218 200826 2454
rect 201062 2218 201146 2454
rect 201382 2218 201414 2454
rect 200794 2134 201414 2218
rect 200794 1898 200826 2134
rect 201062 1898 201146 2134
rect 201382 1898 201414 2134
rect 200794 -346 201414 1898
rect 200794 -582 200826 -346
rect 201062 -582 201146 -346
rect 201382 -582 201414 -346
rect 200794 -666 201414 -582
rect 200794 -902 200826 -666
rect 201062 -902 201146 -666
rect 201382 -902 201414 -666
rect 200794 -1894 201414 -902
rect 204514 686174 205134 706202
rect 204514 685938 204546 686174
rect 204782 685938 204866 686174
rect 205102 685938 205134 686174
rect 204514 685854 205134 685938
rect 204514 685618 204546 685854
rect 204782 685618 204866 685854
rect 205102 685618 205134 685854
rect 204514 646174 205134 685618
rect 204514 645938 204546 646174
rect 204782 645938 204866 646174
rect 205102 645938 205134 646174
rect 204514 645854 205134 645938
rect 204514 645618 204546 645854
rect 204782 645618 204866 645854
rect 205102 645618 205134 645854
rect 204514 606174 205134 645618
rect 204514 605938 204546 606174
rect 204782 605938 204866 606174
rect 205102 605938 205134 606174
rect 204514 605854 205134 605938
rect 204514 605618 204546 605854
rect 204782 605618 204866 605854
rect 205102 605618 205134 605854
rect 204514 566174 205134 605618
rect 204514 565938 204546 566174
rect 204782 565938 204866 566174
rect 205102 565938 205134 566174
rect 204514 565854 205134 565938
rect 204514 565618 204546 565854
rect 204782 565618 204866 565854
rect 205102 565618 205134 565854
rect 204514 526174 205134 565618
rect 204514 525938 204546 526174
rect 204782 525938 204866 526174
rect 205102 525938 205134 526174
rect 204514 525854 205134 525938
rect 204514 525618 204546 525854
rect 204782 525618 204866 525854
rect 205102 525618 205134 525854
rect 204514 486174 205134 525618
rect 204514 485938 204546 486174
rect 204782 485938 204866 486174
rect 205102 485938 205134 486174
rect 204514 485854 205134 485938
rect 204514 485618 204546 485854
rect 204782 485618 204866 485854
rect 205102 485618 205134 485854
rect 204514 446174 205134 485618
rect 204514 445938 204546 446174
rect 204782 445938 204866 446174
rect 205102 445938 205134 446174
rect 204514 445854 205134 445938
rect 204514 445618 204546 445854
rect 204782 445618 204866 445854
rect 205102 445618 205134 445854
rect 204514 406174 205134 445618
rect 204514 405938 204546 406174
rect 204782 405938 204866 406174
rect 205102 405938 205134 406174
rect 204514 405854 205134 405938
rect 204514 405618 204546 405854
rect 204782 405618 204866 405854
rect 205102 405618 205134 405854
rect 204514 366174 205134 405618
rect 204514 365938 204546 366174
rect 204782 365938 204866 366174
rect 205102 365938 205134 366174
rect 204514 365854 205134 365938
rect 204514 365618 204546 365854
rect 204782 365618 204866 365854
rect 205102 365618 205134 365854
rect 204514 326174 205134 365618
rect 204514 325938 204546 326174
rect 204782 325938 204866 326174
rect 205102 325938 205134 326174
rect 204514 325854 205134 325938
rect 204514 325618 204546 325854
rect 204782 325618 204866 325854
rect 205102 325618 205134 325854
rect 204514 286174 205134 325618
rect 204514 285938 204546 286174
rect 204782 285938 204866 286174
rect 205102 285938 205134 286174
rect 204514 285854 205134 285938
rect 204514 285618 204546 285854
rect 204782 285618 204866 285854
rect 205102 285618 205134 285854
rect 204514 246174 205134 285618
rect 204514 245938 204546 246174
rect 204782 245938 204866 246174
rect 205102 245938 205134 246174
rect 204514 245854 205134 245938
rect 204514 245618 204546 245854
rect 204782 245618 204866 245854
rect 205102 245618 205134 245854
rect 204514 206174 205134 245618
rect 204514 205938 204546 206174
rect 204782 205938 204866 206174
rect 205102 205938 205134 206174
rect 204514 205854 205134 205938
rect 204514 205618 204546 205854
rect 204782 205618 204866 205854
rect 205102 205618 205134 205854
rect 204514 166174 205134 205618
rect 204514 165938 204546 166174
rect 204782 165938 204866 166174
rect 205102 165938 205134 166174
rect 204514 165854 205134 165938
rect 204514 165618 204546 165854
rect 204782 165618 204866 165854
rect 205102 165618 205134 165854
rect 204514 126174 205134 165618
rect 204514 125938 204546 126174
rect 204782 125938 204866 126174
rect 205102 125938 205134 126174
rect 204514 125854 205134 125938
rect 204514 125618 204546 125854
rect 204782 125618 204866 125854
rect 205102 125618 205134 125854
rect 204514 86174 205134 125618
rect 204514 85938 204546 86174
rect 204782 85938 204866 86174
rect 205102 85938 205134 86174
rect 204514 85854 205134 85938
rect 204514 85618 204546 85854
rect 204782 85618 204866 85854
rect 205102 85618 205134 85854
rect 204514 46174 205134 85618
rect 204514 45938 204546 46174
rect 204782 45938 204866 46174
rect 205102 45938 205134 46174
rect 204514 45854 205134 45938
rect 204514 45618 204546 45854
rect 204782 45618 204866 45854
rect 205102 45618 205134 45854
rect 204514 6174 205134 45618
rect 204514 5938 204546 6174
rect 204782 5938 204866 6174
rect 205102 5938 205134 6174
rect 204514 5854 205134 5938
rect 204514 5618 204546 5854
rect 204782 5618 204866 5854
rect 205102 5618 205134 5854
rect 204514 -2266 205134 5618
rect 204514 -2502 204546 -2266
rect 204782 -2502 204866 -2266
rect 205102 -2502 205134 -2266
rect 204514 -2586 205134 -2502
rect 204514 -2822 204546 -2586
rect 204782 -2822 204866 -2586
rect 205102 -2822 205134 -2586
rect 204514 -3814 205134 -2822
rect 208234 689894 208854 708122
rect 208234 689658 208266 689894
rect 208502 689658 208586 689894
rect 208822 689658 208854 689894
rect 208234 689574 208854 689658
rect 208234 689338 208266 689574
rect 208502 689338 208586 689574
rect 208822 689338 208854 689574
rect 208234 649894 208854 689338
rect 208234 649658 208266 649894
rect 208502 649658 208586 649894
rect 208822 649658 208854 649894
rect 208234 649574 208854 649658
rect 208234 649338 208266 649574
rect 208502 649338 208586 649574
rect 208822 649338 208854 649574
rect 208234 609894 208854 649338
rect 208234 609658 208266 609894
rect 208502 609658 208586 609894
rect 208822 609658 208854 609894
rect 208234 609574 208854 609658
rect 208234 609338 208266 609574
rect 208502 609338 208586 609574
rect 208822 609338 208854 609574
rect 208234 569894 208854 609338
rect 208234 569658 208266 569894
rect 208502 569658 208586 569894
rect 208822 569658 208854 569894
rect 208234 569574 208854 569658
rect 208234 569338 208266 569574
rect 208502 569338 208586 569574
rect 208822 569338 208854 569574
rect 208234 529894 208854 569338
rect 208234 529658 208266 529894
rect 208502 529658 208586 529894
rect 208822 529658 208854 529894
rect 208234 529574 208854 529658
rect 208234 529338 208266 529574
rect 208502 529338 208586 529574
rect 208822 529338 208854 529574
rect 208234 489894 208854 529338
rect 208234 489658 208266 489894
rect 208502 489658 208586 489894
rect 208822 489658 208854 489894
rect 208234 489574 208854 489658
rect 208234 489338 208266 489574
rect 208502 489338 208586 489574
rect 208822 489338 208854 489574
rect 208234 449894 208854 489338
rect 208234 449658 208266 449894
rect 208502 449658 208586 449894
rect 208822 449658 208854 449894
rect 208234 449574 208854 449658
rect 208234 449338 208266 449574
rect 208502 449338 208586 449574
rect 208822 449338 208854 449574
rect 208234 409894 208854 449338
rect 208234 409658 208266 409894
rect 208502 409658 208586 409894
rect 208822 409658 208854 409894
rect 208234 409574 208854 409658
rect 208234 409338 208266 409574
rect 208502 409338 208586 409574
rect 208822 409338 208854 409574
rect 208234 369894 208854 409338
rect 208234 369658 208266 369894
rect 208502 369658 208586 369894
rect 208822 369658 208854 369894
rect 208234 369574 208854 369658
rect 208234 369338 208266 369574
rect 208502 369338 208586 369574
rect 208822 369338 208854 369574
rect 208234 329894 208854 369338
rect 208234 329658 208266 329894
rect 208502 329658 208586 329894
rect 208822 329658 208854 329894
rect 208234 329574 208854 329658
rect 208234 329338 208266 329574
rect 208502 329338 208586 329574
rect 208822 329338 208854 329574
rect 208234 289894 208854 329338
rect 208234 289658 208266 289894
rect 208502 289658 208586 289894
rect 208822 289658 208854 289894
rect 208234 289574 208854 289658
rect 208234 289338 208266 289574
rect 208502 289338 208586 289574
rect 208822 289338 208854 289574
rect 208234 249894 208854 289338
rect 208234 249658 208266 249894
rect 208502 249658 208586 249894
rect 208822 249658 208854 249894
rect 208234 249574 208854 249658
rect 208234 249338 208266 249574
rect 208502 249338 208586 249574
rect 208822 249338 208854 249574
rect 208234 209894 208854 249338
rect 208234 209658 208266 209894
rect 208502 209658 208586 209894
rect 208822 209658 208854 209894
rect 208234 209574 208854 209658
rect 208234 209338 208266 209574
rect 208502 209338 208586 209574
rect 208822 209338 208854 209574
rect 208234 169894 208854 209338
rect 208234 169658 208266 169894
rect 208502 169658 208586 169894
rect 208822 169658 208854 169894
rect 208234 169574 208854 169658
rect 208234 169338 208266 169574
rect 208502 169338 208586 169574
rect 208822 169338 208854 169574
rect 208234 129894 208854 169338
rect 208234 129658 208266 129894
rect 208502 129658 208586 129894
rect 208822 129658 208854 129894
rect 208234 129574 208854 129658
rect 208234 129338 208266 129574
rect 208502 129338 208586 129574
rect 208822 129338 208854 129574
rect 208234 89894 208854 129338
rect 208234 89658 208266 89894
rect 208502 89658 208586 89894
rect 208822 89658 208854 89894
rect 208234 89574 208854 89658
rect 208234 89338 208266 89574
rect 208502 89338 208586 89574
rect 208822 89338 208854 89574
rect 208234 49894 208854 89338
rect 208234 49658 208266 49894
rect 208502 49658 208586 49894
rect 208822 49658 208854 49894
rect 208234 49574 208854 49658
rect 208234 49338 208266 49574
rect 208502 49338 208586 49574
rect 208822 49338 208854 49574
rect 208234 9894 208854 49338
rect 208234 9658 208266 9894
rect 208502 9658 208586 9894
rect 208822 9658 208854 9894
rect 208234 9574 208854 9658
rect 208234 9338 208266 9574
rect 208502 9338 208586 9574
rect 208822 9338 208854 9574
rect 208234 -4186 208854 9338
rect 208234 -4422 208266 -4186
rect 208502 -4422 208586 -4186
rect 208822 -4422 208854 -4186
rect 208234 -4506 208854 -4422
rect 208234 -4742 208266 -4506
rect 208502 -4742 208586 -4506
rect 208822 -4742 208854 -4506
rect 208234 -5734 208854 -4742
rect 211954 693614 212574 710042
rect 231954 711558 232574 711590
rect 231954 711322 231986 711558
rect 232222 711322 232306 711558
rect 232542 711322 232574 711558
rect 231954 711238 232574 711322
rect 231954 711002 231986 711238
rect 232222 711002 232306 711238
rect 232542 711002 232574 711238
rect 228234 709638 228854 709670
rect 228234 709402 228266 709638
rect 228502 709402 228586 709638
rect 228822 709402 228854 709638
rect 228234 709318 228854 709402
rect 228234 709082 228266 709318
rect 228502 709082 228586 709318
rect 228822 709082 228854 709318
rect 224514 707718 225134 707750
rect 224514 707482 224546 707718
rect 224782 707482 224866 707718
rect 225102 707482 225134 707718
rect 224514 707398 225134 707482
rect 224514 707162 224546 707398
rect 224782 707162 224866 707398
rect 225102 707162 225134 707398
rect 211954 693378 211986 693614
rect 212222 693378 212306 693614
rect 212542 693378 212574 693614
rect 211954 693294 212574 693378
rect 211954 693058 211986 693294
rect 212222 693058 212306 693294
rect 212542 693058 212574 693294
rect 211954 653614 212574 693058
rect 211954 653378 211986 653614
rect 212222 653378 212306 653614
rect 212542 653378 212574 653614
rect 211954 653294 212574 653378
rect 211954 653058 211986 653294
rect 212222 653058 212306 653294
rect 212542 653058 212574 653294
rect 211954 613614 212574 653058
rect 211954 613378 211986 613614
rect 212222 613378 212306 613614
rect 212542 613378 212574 613614
rect 211954 613294 212574 613378
rect 211954 613058 211986 613294
rect 212222 613058 212306 613294
rect 212542 613058 212574 613294
rect 211954 573614 212574 613058
rect 211954 573378 211986 573614
rect 212222 573378 212306 573614
rect 212542 573378 212574 573614
rect 211954 573294 212574 573378
rect 211954 573058 211986 573294
rect 212222 573058 212306 573294
rect 212542 573058 212574 573294
rect 211954 533614 212574 573058
rect 211954 533378 211986 533614
rect 212222 533378 212306 533614
rect 212542 533378 212574 533614
rect 211954 533294 212574 533378
rect 211954 533058 211986 533294
rect 212222 533058 212306 533294
rect 212542 533058 212574 533294
rect 211954 493614 212574 533058
rect 211954 493378 211986 493614
rect 212222 493378 212306 493614
rect 212542 493378 212574 493614
rect 211954 493294 212574 493378
rect 211954 493058 211986 493294
rect 212222 493058 212306 493294
rect 212542 493058 212574 493294
rect 211954 453614 212574 493058
rect 211954 453378 211986 453614
rect 212222 453378 212306 453614
rect 212542 453378 212574 453614
rect 211954 453294 212574 453378
rect 211954 453058 211986 453294
rect 212222 453058 212306 453294
rect 212542 453058 212574 453294
rect 211954 413614 212574 453058
rect 211954 413378 211986 413614
rect 212222 413378 212306 413614
rect 212542 413378 212574 413614
rect 211954 413294 212574 413378
rect 211954 413058 211986 413294
rect 212222 413058 212306 413294
rect 212542 413058 212574 413294
rect 211954 373614 212574 413058
rect 211954 373378 211986 373614
rect 212222 373378 212306 373614
rect 212542 373378 212574 373614
rect 211954 373294 212574 373378
rect 211954 373058 211986 373294
rect 212222 373058 212306 373294
rect 212542 373058 212574 373294
rect 211954 333614 212574 373058
rect 211954 333378 211986 333614
rect 212222 333378 212306 333614
rect 212542 333378 212574 333614
rect 211954 333294 212574 333378
rect 211954 333058 211986 333294
rect 212222 333058 212306 333294
rect 212542 333058 212574 333294
rect 211954 293614 212574 333058
rect 211954 293378 211986 293614
rect 212222 293378 212306 293614
rect 212542 293378 212574 293614
rect 211954 293294 212574 293378
rect 211954 293058 211986 293294
rect 212222 293058 212306 293294
rect 212542 293058 212574 293294
rect 211954 253614 212574 293058
rect 211954 253378 211986 253614
rect 212222 253378 212306 253614
rect 212542 253378 212574 253614
rect 211954 253294 212574 253378
rect 211954 253058 211986 253294
rect 212222 253058 212306 253294
rect 212542 253058 212574 253294
rect 211954 213614 212574 253058
rect 211954 213378 211986 213614
rect 212222 213378 212306 213614
rect 212542 213378 212574 213614
rect 211954 213294 212574 213378
rect 211954 213058 211986 213294
rect 212222 213058 212306 213294
rect 212542 213058 212574 213294
rect 211954 173614 212574 213058
rect 211954 173378 211986 173614
rect 212222 173378 212306 173614
rect 212542 173378 212574 173614
rect 211954 173294 212574 173378
rect 211954 173058 211986 173294
rect 212222 173058 212306 173294
rect 212542 173058 212574 173294
rect 211954 133614 212574 173058
rect 211954 133378 211986 133614
rect 212222 133378 212306 133614
rect 212542 133378 212574 133614
rect 211954 133294 212574 133378
rect 211954 133058 211986 133294
rect 212222 133058 212306 133294
rect 212542 133058 212574 133294
rect 211954 93614 212574 133058
rect 211954 93378 211986 93614
rect 212222 93378 212306 93614
rect 212542 93378 212574 93614
rect 211954 93294 212574 93378
rect 211954 93058 211986 93294
rect 212222 93058 212306 93294
rect 212542 93058 212574 93294
rect 211954 53614 212574 93058
rect 211954 53378 211986 53614
rect 212222 53378 212306 53614
rect 212542 53378 212574 53614
rect 211954 53294 212574 53378
rect 211954 53058 211986 53294
rect 212222 53058 212306 53294
rect 212542 53058 212574 53294
rect 211954 13614 212574 53058
rect 211954 13378 211986 13614
rect 212222 13378 212306 13614
rect 212542 13378 212574 13614
rect 211954 13294 212574 13378
rect 211954 13058 211986 13294
rect 212222 13058 212306 13294
rect 212542 13058 212574 13294
rect 191954 -7302 191986 -7066
rect 192222 -7302 192306 -7066
rect 192542 -7302 192574 -7066
rect 191954 -7386 192574 -7302
rect 191954 -7622 191986 -7386
rect 192222 -7622 192306 -7386
rect 192542 -7622 192574 -7386
rect 191954 -7654 192574 -7622
rect 211954 -6106 212574 13058
rect 220794 705798 221414 705830
rect 220794 705562 220826 705798
rect 221062 705562 221146 705798
rect 221382 705562 221414 705798
rect 220794 705478 221414 705562
rect 220794 705242 220826 705478
rect 221062 705242 221146 705478
rect 221382 705242 221414 705478
rect 220794 662454 221414 705242
rect 220794 662218 220826 662454
rect 221062 662218 221146 662454
rect 221382 662218 221414 662454
rect 220794 662134 221414 662218
rect 220794 661898 220826 662134
rect 221062 661898 221146 662134
rect 221382 661898 221414 662134
rect 220794 622454 221414 661898
rect 220794 622218 220826 622454
rect 221062 622218 221146 622454
rect 221382 622218 221414 622454
rect 220794 622134 221414 622218
rect 220794 621898 220826 622134
rect 221062 621898 221146 622134
rect 221382 621898 221414 622134
rect 220794 582454 221414 621898
rect 220794 582218 220826 582454
rect 221062 582218 221146 582454
rect 221382 582218 221414 582454
rect 220794 582134 221414 582218
rect 220794 581898 220826 582134
rect 221062 581898 221146 582134
rect 221382 581898 221414 582134
rect 220794 542454 221414 581898
rect 220794 542218 220826 542454
rect 221062 542218 221146 542454
rect 221382 542218 221414 542454
rect 220794 542134 221414 542218
rect 220794 541898 220826 542134
rect 221062 541898 221146 542134
rect 221382 541898 221414 542134
rect 220794 502454 221414 541898
rect 220794 502218 220826 502454
rect 221062 502218 221146 502454
rect 221382 502218 221414 502454
rect 220794 502134 221414 502218
rect 220794 501898 220826 502134
rect 221062 501898 221146 502134
rect 221382 501898 221414 502134
rect 220794 462454 221414 501898
rect 220794 462218 220826 462454
rect 221062 462218 221146 462454
rect 221382 462218 221414 462454
rect 220794 462134 221414 462218
rect 220794 461898 220826 462134
rect 221062 461898 221146 462134
rect 221382 461898 221414 462134
rect 220794 422454 221414 461898
rect 220794 422218 220826 422454
rect 221062 422218 221146 422454
rect 221382 422218 221414 422454
rect 220794 422134 221414 422218
rect 220794 421898 220826 422134
rect 221062 421898 221146 422134
rect 221382 421898 221414 422134
rect 220794 382454 221414 421898
rect 220794 382218 220826 382454
rect 221062 382218 221146 382454
rect 221382 382218 221414 382454
rect 220794 382134 221414 382218
rect 220794 381898 220826 382134
rect 221062 381898 221146 382134
rect 221382 381898 221414 382134
rect 220794 342454 221414 381898
rect 220794 342218 220826 342454
rect 221062 342218 221146 342454
rect 221382 342218 221414 342454
rect 220794 342134 221414 342218
rect 220794 341898 220826 342134
rect 221062 341898 221146 342134
rect 221382 341898 221414 342134
rect 220794 302454 221414 341898
rect 220794 302218 220826 302454
rect 221382 302218 221414 302454
rect 220794 302134 221414 302218
rect 220794 301898 220826 302134
rect 221382 301898 221414 302134
rect 220794 262454 221414 301898
rect 220794 262218 220826 262454
rect 221382 262218 221414 262454
rect 220794 262134 221414 262218
rect 220794 261898 220826 262134
rect 221382 261898 221414 262134
rect 220794 222454 221414 261898
rect 220794 222218 220826 222454
rect 221382 222218 221414 222454
rect 220794 222134 221414 222218
rect 220794 221898 220826 222134
rect 221382 221898 221414 222134
rect 220794 182454 221414 221898
rect 220794 182218 220826 182454
rect 221382 182218 221414 182454
rect 220794 182134 221414 182218
rect 220794 181898 220826 182134
rect 221382 181898 221414 182134
rect 220794 142454 221414 181898
rect 220794 142218 220826 142454
rect 221382 142218 221414 142454
rect 220794 142134 221414 142218
rect 220794 141898 220826 142134
rect 221382 141898 221414 142134
rect 220794 102454 221414 141898
rect 220794 102218 220826 102454
rect 221062 102218 221146 102454
rect 221382 102218 221414 102454
rect 220794 102134 221414 102218
rect 220794 101898 220826 102134
rect 221062 101898 221146 102134
rect 221382 101898 221414 102134
rect 220794 62454 221414 101898
rect 220794 62218 220826 62454
rect 221062 62218 221146 62454
rect 221382 62218 221414 62454
rect 220794 62134 221414 62218
rect 220794 61898 220826 62134
rect 221062 61898 221146 62134
rect 221382 61898 221414 62134
rect 220794 22454 221414 61898
rect 220794 22218 220826 22454
rect 221062 22218 221146 22454
rect 221382 22218 221414 22454
rect 220794 22134 221414 22218
rect 220794 21898 220826 22134
rect 221062 21898 221146 22134
rect 221382 21898 221414 22134
rect 220794 -1306 221414 21898
rect 220794 -1542 220826 -1306
rect 221062 -1542 221146 -1306
rect 221382 -1542 221414 -1306
rect 220794 -1626 221414 -1542
rect 220794 -1862 220826 -1626
rect 221062 -1862 221146 -1626
rect 221382 -1862 221414 -1626
rect 220794 -1894 221414 -1862
rect 224514 666174 225134 707162
rect 224514 665938 224546 666174
rect 224782 665938 224866 666174
rect 225102 665938 225134 666174
rect 224514 665854 225134 665938
rect 224514 665618 224546 665854
rect 224782 665618 224866 665854
rect 225102 665618 225134 665854
rect 224514 626174 225134 665618
rect 224514 625938 224546 626174
rect 224782 625938 224866 626174
rect 225102 625938 225134 626174
rect 224514 625854 225134 625938
rect 224514 625618 224546 625854
rect 224782 625618 224866 625854
rect 225102 625618 225134 625854
rect 224514 586174 225134 625618
rect 224514 585938 224546 586174
rect 224782 585938 224866 586174
rect 225102 585938 225134 586174
rect 224514 585854 225134 585938
rect 224514 585618 224546 585854
rect 224782 585618 224866 585854
rect 225102 585618 225134 585854
rect 224514 546174 225134 585618
rect 224514 545938 224546 546174
rect 224782 545938 224866 546174
rect 225102 545938 225134 546174
rect 224514 545854 225134 545938
rect 224514 545618 224546 545854
rect 224782 545618 224866 545854
rect 225102 545618 225134 545854
rect 224514 506174 225134 545618
rect 224514 505938 224546 506174
rect 224782 505938 224866 506174
rect 225102 505938 225134 506174
rect 224514 505854 225134 505938
rect 224514 505618 224546 505854
rect 224782 505618 224866 505854
rect 225102 505618 225134 505854
rect 224514 466174 225134 505618
rect 224514 465938 224546 466174
rect 224782 465938 224866 466174
rect 225102 465938 225134 466174
rect 224514 465854 225134 465938
rect 224514 465618 224546 465854
rect 224782 465618 224866 465854
rect 225102 465618 225134 465854
rect 224514 426174 225134 465618
rect 224514 425938 224546 426174
rect 224782 425938 224866 426174
rect 225102 425938 225134 426174
rect 224514 425854 225134 425938
rect 224514 425618 224546 425854
rect 224782 425618 224866 425854
rect 225102 425618 225134 425854
rect 224514 386174 225134 425618
rect 224514 385938 224546 386174
rect 224782 385938 224866 386174
rect 225102 385938 225134 386174
rect 224514 385854 225134 385938
rect 224514 385618 224546 385854
rect 224782 385618 224866 385854
rect 225102 385618 225134 385854
rect 224514 346174 225134 385618
rect 224514 345938 224546 346174
rect 224782 345938 224866 346174
rect 225102 345938 225134 346174
rect 224514 345854 225134 345938
rect 224514 345618 224546 345854
rect 224782 345618 224866 345854
rect 225102 345618 225134 345854
rect 224514 306174 225134 345618
rect 224514 305938 224546 306174
rect 224782 305938 224866 306174
rect 225102 305938 225134 306174
rect 224514 305854 225134 305938
rect 224514 305618 224546 305854
rect 224782 305618 224866 305854
rect 225102 305618 225134 305854
rect 224514 266174 225134 305618
rect 224514 265938 224546 266174
rect 224782 265938 224866 266174
rect 225102 265938 225134 266174
rect 224514 265854 225134 265938
rect 224514 265618 224546 265854
rect 224782 265618 224866 265854
rect 225102 265618 225134 265854
rect 224514 226174 225134 265618
rect 224514 225938 224546 226174
rect 224782 225938 224866 226174
rect 225102 225938 225134 226174
rect 224514 225854 225134 225938
rect 224514 225618 224546 225854
rect 224782 225618 224866 225854
rect 225102 225618 225134 225854
rect 224514 186174 225134 225618
rect 224514 185938 224546 186174
rect 224782 185938 224866 186174
rect 225102 185938 225134 186174
rect 224514 185854 225134 185938
rect 224514 185618 224546 185854
rect 224782 185618 224866 185854
rect 225102 185618 225134 185854
rect 224514 146174 225134 185618
rect 224514 145938 224546 146174
rect 224782 145938 224866 146174
rect 225102 145938 225134 146174
rect 224514 145854 225134 145938
rect 224514 145618 224546 145854
rect 224782 145618 224866 145854
rect 225102 145618 225134 145854
rect 224514 106174 225134 145618
rect 224514 105938 224546 106174
rect 224782 105938 224866 106174
rect 225102 105938 225134 106174
rect 224514 105854 225134 105938
rect 224514 105618 224546 105854
rect 224782 105618 224866 105854
rect 225102 105618 225134 105854
rect 224514 66174 225134 105618
rect 224514 65938 224546 66174
rect 224782 65938 224866 66174
rect 225102 65938 225134 66174
rect 224514 65854 225134 65938
rect 224514 65618 224546 65854
rect 224782 65618 224866 65854
rect 225102 65618 225134 65854
rect 224514 26174 225134 65618
rect 224514 25938 224546 26174
rect 224782 25938 224866 26174
rect 225102 25938 225134 26174
rect 224514 25854 225134 25938
rect 224514 25618 224546 25854
rect 224782 25618 224866 25854
rect 225102 25618 225134 25854
rect 224514 -3226 225134 25618
rect 224514 -3462 224546 -3226
rect 224782 -3462 224866 -3226
rect 225102 -3462 225134 -3226
rect 224514 -3546 225134 -3462
rect 224514 -3782 224546 -3546
rect 224782 -3782 224866 -3546
rect 225102 -3782 225134 -3546
rect 224514 -3814 225134 -3782
rect 228234 669894 228854 709082
rect 228234 669658 228266 669894
rect 228502 669658 228586 669894
rect 228822 669658 228854 669894
rect 228234 669574 228854 669658
rect 228234 669338 228266 669574
rect 228502 669338 228586 669574
rect 228822 669338 228854 669574
rect 228234 629894 228854 669338
rect 228234 629658 228266 629894
rect 228502 629658 228586 629894
rect 228822 629658 228854 629894
rect 228234 629574 228854 629658
rect 228234 629338 228266 629574
rect 228502 629338 228586 629574
rect 228822 629338 228854 629574
rect 228234 589894 228854 629338
rect 228234 589658 228266 589894
rect 228502 589658 228586 589894
rect 228822 589658 228854 589894
rect 228234 589574 228854 589658
rect 228234 589338 228266 589574
rect 228502 589338 228586 589574
rect 228822 589338 228854 589574
rect 228234 549894 228854 589338
rect 228234 549658 228266 549894
rect 228502 549658 228586 549894
rect 228822 549658 228854 549894
rect 228234 549574 228854 549658
rect 228234 549338 228266 549574
rect 228502 549338 228586 549574
rect 228822 549338 228854 549574
rect 228234 509894 228854 549338
rect 228234 509658 228266 509894
rect 228502 509658 228586 509894
rect 228822 509658 228854 509894
rect 228234 509574 228854 509658
rect 228234 509338 228266 509574
rect 228502 509338 228586 509574
rect 228822 509338 228854 509574
rect 228234 469894 228854 509338
rect 228234 469658 228266 469894
rect 228502 469658 228586 469894
rect 228822 469658 228854 469894
rect 228234 469574 228854 469658
rect 228234 469338 228266 469574
rect 228502 469338 228586 469574
rect 228822 469338 228854 469574
rect 228234 429894 228854 469338
rect 228234 429658 228266 429894
rect 228502 429658 228586 429894
rect 228822 429658 228854 429894
rect 228234 429574 228854 429658
rect 228234 429338 228266 429574
rect 228502 429338 228586 429574
rect 228822 429338 228854 429574
rect 228234 389894 228854 429338
rect 228234 389658 228266 389894
rect 228502 389658 228586 389894
rect 228822 389658 228854 389894
rect 228234 389574 228854 389658
rect 228234 389338 228266 389574
rect 228502 389338 228586 389574
rect 228822 389338 228854 389574
rect 228234 349894 228854 389338
rect 228234 349658 228266 349894
rect 228502 349658 228586 349894
rect 228822 349658 228854 349894
rect 228234 349574 228854 349658
rect 228234 349338 228266 349574
rect 228502 349338 228586 349574
rect 228822 349338 228854 349574
rect 228234 309894 228854 349338
rect 228234 309658 228266 309894
rect 228502 309658 228586 309894
rect 228822 309658 228854 309894
rect 228234 309574 228854 309658
rect 228234 309338 228266 309574
rect 228502 309338 228586 309574
rect 228822 309338 228854 309574
rect 228234 269894 228854 309338
rect 228234 269658 228266 269894
rect 228502 269658 228586 269894
rect 228822 269658 228854 269894
rect 228234 269574 228854 269658
rect 228234 269338 228266 269574
rect 228502 269338 228586 269574
rect 228822 269338 228854 269574
rect 228234 229894 228854 269338
rect 228234 229658 228266 229894
rect 228502 229658 228586 229894
rect 228822 229658 228854 229894
rect 228234 229574 228854 229658
rect 228234 229338 228266 229574
rect 228502 229338 228586 229574
rect 228822 229338 228854 229574
rect 228234 189894 228854 229338
rect 228234 189658 228266 189894
rect 228502 189658 228586 189894
rect 228822 189658 228854 189894
rect 228234 189574 228854 189658
rect 228234 189338 228266 189574
rect 228502 189338 228586 189574
rect 228822 189338 228854 189574
rect 228234 149894 228854 189338
rect 228234 149658 228266 149894
rect 228502 149658 228586 149894
rect 228822 149658 228854 149894
rect 228234 149574 228854 149658
rect 228234 149338 228266 149574
rect 228502 149338 228586 149574
rect 228822 149338 228854 149574
rect 228234 109894 228854 149338
rect 228234 109658 228266 109894
rect 228502 109658 228586 109894
rect 228822 109658 228854 109894
rect 228234 109574 228854 109658
rect 228234 109338 228266 109574
rect 228502 109338 228586 109574
rect 228822 109338 228854 109574
rect 228234 69894 228854 109338
rect 228234 69658 228266 69894
rect 228502 69658 228586 69894
rect 228822 69658 228854 69894
rect 228234 69574 228854 69658
rect 228234 69338 228266 69574
rect 228502 69338 228586 69574
rect 228822 69338 228854 69574
rect 228234 29894 228854 69338
rect 228234 29658 228266 29894
rect 228502 29658 228586 29894
rect 228822 29658 228854 29894
rect 228234 29574 228854 29658
rect 228234 29338 228266 29574
rect 228502 29338 228586 29574
rect 228822 29338 228854 29574
rect 228234 -5146 228854 29338
rect 228234 -5382 228266 -5146
rect 228502 -5382 228586 -5146
rect 228822 -5382 228854 -5146
rect 228234 -5466 228854 -5382
rect 228234 -5702 228266 -5466
rect 228502 -5702 228586 -5466
rect 228822 -5702 228854 -5466
rect 228234 -5734 228854 -5702
rect 231954 673614 232574 711002
rect 251954 710598 252574 711590
rect 251954 710362 251986 710598
rect 252222 710362 252306 710598
rect 252542 710362 252574 710598
rect 251954 710278 252574 710362
rect 251954 710042 251986 710278
rect 252222 710042 252306 710278
rect 252542 710042 252574 710278
rect 248234 708678 248854 709670
rect 248234 708442 248266 708678
rect 248502 708442 248586 708678
rect 248822 708442 248854 708678
rect 248234 708358 248854 708442
rect 248234 708122 248266 708358
rect 248502 708122 248586 708358
rect 248822 708122 248854 708358
rect 244514 706758 245134 707750
rect 244514 706522 244546 706758
rect 244782 706522 244866 706758
rect 245102 706522 245134 706758
rect 244514 706438 245134 706522
rect 244514 706202 244546 706438
rect 244782 706202 244866 706438
rect 245102 706202 245134 706438
rect 231954 673378 231986 673614
rect 232222 673378 232306 673614
rect 232542 673378 232574 673614
rect 231954 673294 232574 673378
rect 231954 673058 231986 673294
rect 232222 673058 232306 673294
rect 232542 673058 232574 673294
rect 231954 633614 232574 673058
rect 231954 633378 231986 633614
rect 232222 633378 232306 633614
rect 232542 633378 232574 633614
rect 231954 633294 232574 633378
rect 231954 633058 231986 633294
rect 232222 633058 232306 633294
rect 232542 633058 232574 633294
rect 231954 593614 232574 633058
rect 231954 593378 231986 593614
rect 232222 593378 232306 593614
rect 232542 593378 232574 593614
rect 231954 593294 232574 593378
rect 231954 593058 231986 593294
rect 232222 593058 232306 593294
rect 232542 593058 232574 593294
rect 231954 553614 232574 593058
rect 231954 553378 231986 553614
rect 232222 553378 232306 553614
rect 232542 553378 232574 553614
rect 231954 553294 232574 553378
rect 231954 553058 231986 553294
rect 232222 553058 232306 553294
rect 232542 553058 232574 553294
rect 231954 513614 232574 553058
rect 231954 513378 231986 513614
rect 232222 513378 232306 513614
rect 232542 513378 232574 513614
rect 231954 513294 232574 513378
rect 231954 513058 231986 513294
rect 232222 513058 232306 513294
rect 232542 513058 232574 513294
rect 231954 473614 232574 513058
rect 231954 473378 231986 473614
rect 232222 473378 232306 473614
rect 232542 473378 232574 473614
rect 231954 473294 232574 473378
rect 231954 473058 231986 473294
rect 232222 473058 232306 473294
rect 232542 473058 232574 473294
rect 231954 433614 232574 473058
rect 231954 433378 231986 433614
rect 232222 433378 232306 433614
rect 232542 433378 232574 433614
rect 231954 433294 232574 433378
rect 231954 433058 231986 433294
rect 232222 433058 232306 433294
rect 232542 433058 232574 433294
rect 231954 393614 232574 433058
rect 231954 393378 231986 393614
rect 232222 393378 232306 393614
rect 232542 393378 232574 393614
rect 231954 393294 232574 393378
rect 231954 393058 231986 393294
rect 232222 393058 232306 393294
rect 232542 393058 232574 393294
rect 231954 353614 232574 393058
rect 231954 353378 231986 353614
rect 232222 353378 232306 353614
rect 232542 353378 232574 353614
rect 231954 353294 232574 353378
rect 231954 353058 231986 353294
rect 232222 353058 232306 353294
rect 232542 353058 232574 353294
rect 231954 313614 232574 353058
rect 240794 704838 241414 705830
rect 240794 704602 240826 704838
rect 241062 704602 241146 704838
rect 241382 704602 241414 704838
rect 240794 704518 241414 704602
rect 240794 704282 240826 704518
rect 241062 704282 241146 704518
rect 241382 704282 241414 704518
rect 240794 682454 241414 704282
rect 240794 682218 240826 682454
rect 241062 682218 241146 682454
rect 241382 682218 241414 682454
rect 240794 682134 241414 682218
rect 240794 681898 240826 682134
rect 241062 681898 241146 682134
rect 241382 681898 241414 682134
rect 240794 642454 241414 681898
rect 240794 642218 240826 642454
rect 241062 642218 241146 642454
rect 241382 642218 241414 642454
rect 240794 642134 241414 642218
rect 240794 641898 240826 642134
rect 241062 641898 241146 642134
rect 241382 641898 241414 642134
rect 240794 602454 241414 641898
rect 240794 602218 240826 602454
rect 241062 602218 241146 602454
rect 241382 602218 241414 602454
rect 240794 602134 241414 602218
rect 240794 601898 240826 602134
rect 241062 601898 241146 602134
rect 241382 601898 241414 602134
rect 240794 562454 241414 601898
rect 240794 562218 240826 562454
rect 241062 562218 241146 562454
rect 241382 562218 241414 562454
rect 240794 562134 241414 562218
rect 240794 561898 240826 562134
rect 241062 561898 241146 562134
rect 241382 561898 241414 562134
rect 240794 522454 241414 561898
rect 240794 522218 240826 522454
rect 241062 522218 241146 522454
rect 241382 522218 241414 522454
rect 240794 522134 241414 522218
rect 240794 521898 240826 522134
rect 241062 521898 241146 522134
rect 241382 521898 241414 522134
rect 240794 482454 241414 521898
rect 240794 482218 240826 482454
rect 241062 482218 241146 482454
rect 241382 482218 241414 482454
rect 240794 482134 241414 482218
rect 240794 481898 240826 482134
rect 241062 481898 241146 482134
rect 241382 481898 241414 482134
rect 240794 442454 241414 481898
rect 240794 442218 240826 442454
rect 241062 442218 241146 442454
rect 241382 442218 241414 442454
rect 240794 442134 241414 442218
rect 240794 441898 240826 442134
rect 241062 441898 241146 442134
rect 241382 441898 241414 442134
rect 240794 402454 241414 441898
rect 240794 402218 240826 402454
rect 241062 402218 241146 402454
rect 241382 402218 241414 402454
rect 240794 402134 241414 402218
rect 240794 401898 240826 402134
rect 241062 401898 241146 402134
rect 241382 401898 241414 402134
rect 240794 362454 241414 401898
rect 240794 362218 240826 362454
rect 241062 362218 241146 362454
rect 241382 362218 241414 362454
rect 240794 362134 241414 362218
rect 240794 361898 240826 362134
rect 241062 361898 241146 362134
rect 241382 361898 241414 362134
rect 240794 322454 241414 361898
rect 240794 322218 240826 322454
rect 241062 322218 241146 322454
rect 241382 322218 241414 322454
rect 240794 322134 241414 322218
rect 240794 321898 240826 322134
rect 241062 321898 241146 322134
rect 241382 321898 241414 322134
rect 232819 319428 232885 319429
rect 232819 319364 232820 319428
rect 232884 319364 232885 319428
rect 232819 319363 232885 319364
rect 231954 313378 231986 313614
rect 232222 313378 232306 313614
rect 232542 313378 232574 313614
rect 231954 313294 232574 313378
rect 231954 313058 231986 313294
rect 232222 313058 232306 313294
rect 232542 313058 232574 313294
rect 231954 273614 232574 313058
rect 231954 273378 231986 273614
rect 232222 273378 232306 273614
rect 232542 273378 232574 273614
rect 231954 273294 232574 273378
rect 231954 273058 231986 273294
rect 232222 273058 232306 273294
rect 232542 273058 232574 273294
rect 231954 233614 232574 273058
rect 231954 233378 231986 233614
rect 232222 233378 232306 233614
rect 232542 233378 232574 233614
rect 231954 233294 232574 233378
rect 231954 233058 231986 233294
rect 232222 233058 232306 233294
rect 232542 233058 232574 233294
rect 231954 193614 232574 233058
rect 231954 193378 231986 193614
rect 232222 193378 232306 193614
rect 232542 193378 232574 193614
rect 231954 193294 232574 193378
rect 231954 193058 231986 193294
rect 232222 193058 232306 193294
rect 232542 193058 232574 193294
rect 231954 153614 232574 193058
rect 231954 153378 231986 153614
rect 232222 153378 232306 153614
rect 232542 153378 232574 153614
rect 231954 153294 232574 153378
rect 231954 153058 231986 153294
rect 232222 153058 232306 153294
rect 232542 153058 232574 153294
rect 231954 113614 232574 153058
rect 231954 113378 231986 113614
rect 232222 113378 232306 113614
rect 232542 113378 232574 113614
rect 231954 113294 232574 113378
rect 231954 113058 231986 113294
rect 232222 113058 232306 113294
rect 232542 113058 232574 113294
rect 231954 73614 232574 113058
rect 231954 73378 231986 73614
rect 232222 73378 232306 73614
rect 232542 73378 232574 73614
rect 231954 73294 232574 73378
rect 231954 73058 231986 73294
rect 232222 73058 232306 73294
rect 232542 73058 232574 73294
rect 231954 33614 232574 73058
rect 231954 33378 231986 33614
rect 232222 33378 232306 33614
rect 232542 33378 232574 33614
rect 231954 33294 232574 33378
rect 231954 33058 231986 33294
rect 232222 33058 232306 33294
rect 232542 33058 232574 33294
rect 211954 -6342 211986 -6106
rect 212222 -6342 212306 -6106
rect 212542 -6342 212574 -6106
rect 211954 -6426 212574 -6342
rect 211954 -6662 211986 -6426
rect 212222 -6662 212306 -6426
rect 212542 -6662 212574 -6426
rect 211954 -7654 212574 -6662
rect 231954 -7066 232574 33058
rect 232822 3909 232882 319363
rect 240794 282454 241414 321898
rect 240794 282218 240826 282454
rect 241382 282218 241414 282454
rect 240794 282134 241414 282218
rect 240794 281898 240826 282134
rect 241382 281898 241414 282134
rect 240794 242454 241414 281898
rect 240794 242218 240826 242454
rect 241382 242218 241414 242454
rect 240794 242134 241414 242218
rect 240794 241898 240826 242134
rect 241382 241898 241414 242134
rect 240794 202454 241414 241898
rect 240794 202218 240826 202454
rect 241382 202218 241414 202454
rect 240794 202134 241414 202218
rect 240794 201898 240826 202134
rect 241382 201898 241414 202134
rect 240794 162454 241414 201898
rect 240794 162218 240826 162454
rect 241382 162218 241414 162454
rect 240794 162134 241414 162218
rect 240794 161898 240826 162134
rect 241382 161898 241414 162134
rect 240794 122454 241414 161898
rect 240794 122218 240826 122454
rect 241062 122218 241146 122454
rect 241382 122218 241414 122454
rect 240794 122134 241414 122218
rect 240794 121898 240826 122134
rect 241062 121898 241146 122134
rect 241382 121898 241414 122134
rect 240794 82454 241414 121898
rect 240794 82218 240826 82454
rect 241062 82218 241146 82454
rect 241382 82218 241414 82454
rect 240794 82134 241414 82218
rect 240794 81898 240826 82134
rect 241062 81898 241146 82134
rect 241382 81898 241414 82134
rect 240794 42454 241414 81898
rect 240794 42218 240826 42454
rect 241062 42218 241146 42454
rect 241382 42218 241414 42454
rect 240794 42134 241414 42218
rect 240794 41898 240826 42134
rect 241062 41898 241146 42134
rect 241382 41898 241414 42134
rect 232819 3908 232885 3909
rect 232819 3844 232820 3908
rect 232884 3844 232885 3908
rect 232819 3843 232885 3844
rect 240794 2454 241414 41898
rect 240794 2218 240826 2454
rect 241062 2218 241146 2454
rect 241382 2218 241414 2454
rect 240794 2134 241414 2218
rect 240794 1898 240826 2134
rect 241062 1898 241146 2134
rect 241382 1898 241414 2134
rect 240794 -346 241414 1898
rect 240794 -582 240826 -346
rect 241062 -582 241146 -346
rect 241382 -582 241414 -346
rect 240794 -666 241414 -582
rect 240794 -902 240826 -666
rect 241062 -902 241146 -666
rect 241382 -902 241414 -666
rect 240794 -1894 241414 -902
rect 244514 686174 245134 706202
rect 244514 685938 244546 686174
rect 244782 685938 244866 686174
rect 245102 685938 245134 686174
rect 244514 685854 245134 685938
rect 244514 685618 244546 685854
rect 244782 685618 244866 685854
rect 245102 685618 245134 685854
rect 244514 646174 245134 685618
rect 244514 645938 244546 646174
rect 244782 645938 244866 646174
rect 245102 645938 245134 646174
rect 244514 645854 245134 645938
rect 244514 645618 244546 645854
rect 244782 645618 244866 645854
rect 245102 645618 245134 645854
rect 244514 606174 245134 645618
rect 244514 605938 244546 606174
rect 244782 605938 244866 606174
rect 245102 605938 245134 606174
rect 244514 605854 245134 605938
rect 244514 605618 244546 605854
rect 244782 605618 244866 605854
rect 245102 605618 245134 605854
rect 244514 566174 245134 605618
rect 244514 565938 244546 566174
rect 244782 565938 244866 566174
rect 245102 565938 245134 566174
rect 244514 565854 245134 565938
rect 244514 565618 244546 565854
rect 244782 565618 244866 565854
rect 245102 565618 245134 565854
rect 244514 526174 245134 565618
rect 244514 525938 244546 526174
rect 244782 525938 244866 526174
rect 245102 525938 245134 526174
rect 244514 525854 245134 525938
rect 244514 525618 244546 525854
rect 244782 525618 244866 525854
rect 245102 525618 245134 525854
rect 244514 486174 245134 525618
rect 244514 485938 244546 486174
rect 244782 485938 244866 486174
rect 245102 485938 245134 486174
rect 244514 485854 245134 485938
rect 244514 485618 244546 485854
rect 244782 485618 244866 485854
rect 245102 485618 245134 485854
rect 244514 446174 245134 485618
rect 244514 445938 244546 446174
rect 244782 445938 244866 446174
rect 245102 445938 245134 446174
rect 244514 445854 245134 445938
rect 244514 445618 244546 445854
rect 244782 445618 244866 445854
rect 245102 445618 245134 445854
rect 244514 406174 245134 445618
rect 244514 405938 244546 406174
rect 244782 405938 244866 406174
rect 245102 405938 245134 406174
rect 244514 405854 245134 405938
rect 244514 405618 244546 405854
rect 244782 405618 244866 405854
rect 245102 405618 245134 405854
rect 244514 366174 245134 405618
rect 244514 365938 244546 366174
rect 244782 365938 244866 366174
rect 245102 365938 245134 366174
rect 244514 365854 245134 365938
rect 244514 365618 244546 365854
rect 244782 365618 244866 365854
rect 245102 365618 245134 365854
rect 244514 326174 245134 365618
rect 244514 325938 244546 326174
rect 244782 325938 244866 326174
rect 245102 325938 245134 326174
rect 244514 325854 245134 325938
rect 244514 325618 244546 325854
rect 244782 325618 244866 325854
rect 245102 325618 245134 325854
rect 244514 286174 245134 325618
rect 244514 285938 244546 286174
rect 244782 285938 244866 286174
rect 245102 285938 245134 286174
rect 244514 285854 245134 285938
rect 244514 285618 244546 285854
rect 244782 285618 244866 285854
rect 245102 285618 245134 285854
rect 244514 246174 245134 285618
rect 244514 245938 244546 246174
rect 244782 245938 244866 246174
rect 245102 245938 245134 246174
rect 244514 245854 245134 245938
rect 244514 245618 244546 245854
rect 244782 245618 244866 245854
rect 245102 245618 245134 245854
rect 244514 206174 245134 245618
rect 244514 205938 244546 206174
rect 244782 205938 244866 206174
rect 245102 205938 245134 206174
rect 244514 205854 245134 205938
rect 244514 205618 244546 205854
rect 244782 205618 244866 205854
rect 245102 205618 245134 205854
rect 244514 166174 245134 205618
rect 244514 165938 244546 166174
rect 244782 165938 244866 166174
rect 245102 165938 245134 166174
rect 244514 165854 245134 165938
rect 244514 165618 244546 165854
rect 244782 165618 244866 165854
rect 245102 165618 245134 165854
rect 244514 126174 245134 165618
rect 244514 125938 244546 126174
rect 244782 125938 244866 126174
rect 245102 125938 245134 126174
rect 244514 125854 245134 125938
rect 244514 125618 244546 125854
rect 244782 125618 244866 125854
rect 245102 125618 245134 125854
rect 244514 86174 245134 125618
rect 244514 85938 244546 86174
rect 244782 85938 244866 86174
rect 245102 85938 245134 86174
rect 244514 85854 245134 85938
rect 244514 85618 244546 85854
rect 244782 85618 244866 85854
rect 245102 85618 245134 85854
rect 244514 46174 245134 85618
rect 244514 45938 244546 46174
rect 244782 45938 244866 46174
rect 245102 45938 245134 46174
rect 244514 45854 245134 45938
rect 244514 45618 244546 45854
rect 244782 45618 244866 45854
rect 245102 45618 245134 45854
rect 244514 6174 245134 45618
rect 244514 5938 244546 6174
rect 244782 5938 244866 6174
rect 245102 5938 245134 6174
rect 244514 5854 245134 5938
rect 244514 5618 244546 5854
rect 244782 5618 244866 5854
rect 245102 5618 245134 5854
rect 244514 -2266 245134 5618
rect 244514 -2502 244546 -2266
rect 244782 -2502 244866 -2266
rect 245102 -2502 245134 -2266
rect 244514 -2586 245134 -2502
rect 244514 -2822 244546 -2586
rect 244782 -2822 244866 -2586
rect 245102 -2822 245134 -2586
rect 244514 -3814 245134 -2822
rect 248234 689894 248854 708122
rect 248234 689658 248266 689894
rect 248502 689658 248586 689894
rect 248822 689658 248854 689894
rect 248234 689574 248854 689658
rect 248234 689338 248266 689574
rect 248502 689338 248586 689574
rect 248822 689338 248854 689574
rect 248234 649894 248854 689338
rect 248234 649658 248266 649894
rect 248502 649658 248586 649894
rect 248822 649658 248854 649894
rect 248234 649574 248854 649658
rect 248234 649338 248266 649574
rect 248502 649338 248586 649574
rect 248822 649338 248854 649574
rect 248234 609894 248854 649338
rect 248234 609658 248266 609894
rect 248502 609658 248586 609894
rect 248822 609658 248854 609894
rect 248234 609574 248854 609658
rect 248234 609338 248266 609574
rect 248502 609338 248586 609574
rect 248822 609338 248854 609574
rect 248234 569894 248854 609338
rect 248234 569658 248266 569894
rect 248502 569658 248586 569894
rect 248822 569658 248854 569894
rect 248234 569574 248854 569658
rect 248234 569338 248266 569574
rect 248502 569338 248586 569574
rect 248822 569338 248854 569574
rect 248234 529894 248854 569338
rect 248234 529658 248266 529894
rect 248502 529658 248586 529894
rect 248822 529658 248854 529894
rect 248234 529574 248854 529658
rect 248234 529338 248266 529574
rect 248502 529338 248586 529574
rect 248822 529338 248854 529574
rect 248234 489894 248854 529338
rect 248234 489658 248266 489894
rect 248502 489658 248586 489894
rect 248822 489658 248854 489894
rect 248234 489574 248854 489658
rect 248234 489338 248266 489574
rect 248502 489338 248586 489574
rect 248822 489338 248854 489574
rect 248234 449894 248854 489338
rect 248234 449658 248266 449894
rect 248502 449658 248586 449894
rect 248822 449658 248854 449894
rect 248234 449574 248854 449658
rect 248234 449338 248266 449574
rect 248502 449338 248586 449574
rect 248822 449338 248854 449574
rect 248234 409894 248854 449338
rect 248234 409658 248266 409894
rect 248502 409658 248586 409894
rect 248822 409658 248854 409894
rect 248234 409574 248854 409658
rect 248234 409338 248266 409574
rect 248502 409338 248586 409574
rect 248822 409338 248854 409574
rect 248234 369894 248854 409338
rect 248234 369658 248266 369894
rect 248502 369658 248586 369894
rect 248822 369658 248854 369894
rect 248234 369574 248854 369658
rect 248234 369338 248266 369574
rect 248502 369338 248586 369574
rect 248822 369338 248854 369574
rect 248234 329894 248854 369338
rect 248234 329658 248266 329894
rect 248502 329658 248586 329894
rect 248822 329658 248854 329894
rect 248234 329574 248854 329658
rect 248234 329338 248266 329574
rect 248502 329338 248586 329574
rect 248822 329338 248854 329574
rect 248234 289894 248854 329338
rect 248234 289658 248266 289894
rect 248502 289658 248586 289894
rect 248822 289658 248854 289894
rect 248234 289574 248854 289658
rect 248234 289338 248266 289574
rect 248502 289338 248586 289574
rect 248822 289338 248854 289574
rect 248234 249894 248854 289338
rect 248234 249658 248266 249894
rect 248502 249658 248586 249894
rect 248822 249658 248854 249894
rect 248234 249574 248854 249658
rect 248234 249338 248266 249574
rect 248502 249338 248586 249574
rect 248822 249338 248854 249574
rect 248234 209894 248854 249338
rect 248234 209658 248266 209894
rect 248502 209658 248586 209894
rect 248822 209658 248854 209894
rect 248234 209574 248854 209658
rect 248234 209338 248266 209574
rect 248502 209338 248586 209574
rect 248822 209338 248854 209574
rect 248234 169894 248854 209338
rect 248234 169658 248266 169894
rect 248502 169658 248586 169894
rect 248822 169658 248854 169894
rect 248234 169574 248854 169658
rect 248234 169338 248266 169574
rect 248502 169338 248586 169574
rect 248822 169338 248854 169574
rect 248234 129894 248854 169338
rect 248234 129658 248266 129894
rect 248502 129658 248586 129894
rect 248822 129658 248854 129894
rect 248234 129574 248854 129658
rect 248234 129338 248266 129574
rect 248502 129338 248586 129574
rect 248822 129338 248854 129574
rect 248234 89894 248854 129338
rect 248234 89658 248266 89894
rect 248502 89658 248586 89894
rect 248822 89658 248854 89894
rect 248234 89574 248854 89658
rect 248234 89338 248266 89574
rect 248502 89338 248586 89574
rect 248822 89338 248854 89574
rect 248234 49894 248854 89338
rect 248234 49658 248266 49894
rect 248502 49658 248586 49894
rect 248822 49658 248854 49894
rect 248234 49574 248854 49658
rect 248234 49338 248266 49574
rect 248502 49338 248586 49574
rect 248822 49338 248854 49574
rect 248234 9894 248854 49338
rect 248234 9658 248266 9894
rect 248502 9658 248586 9894
rect 248822 9658 248854 9894
rect 248234 9574 248854 9658
rect 248234 9338 248266 9574
rect 248502 9338 248586 9574
rect 248822 9338 248854 9574
rect 248234 -4186 248854 9338
rect 248234 -4422 248266 -4186
rect 248502 -4422 248586 -4186
rect 248822 -4422 248854 -4186
rect 248234 -4506 248854 -4422
rect 248234 -4742 248266 -4506
rect 248502 -4742 248586 -4506
rect 248822 -4742 248854 -4506
rect 248234 -5734 248854 -4742
rect 251954 693614 252574 710042
rect 271954 711558 272574 711590
rect 271954 711322 271986 711558
rect 272222 711322 272306 711558
rect 272542 711322 272574 711558
rect 271954 711238 272574 711322
rect 271954 711002 271986 711238
rect 272222 711002 272306 711238
rect 272542 711002 272574 711238
rect 268234 709638 268854 709670
rect 268234 709402 268266 709638
rect 268502 709402 268586 709638
rect 268822 709402 268854 709638
rect 268234 709318 268854 709402
rect 268234 709082 268266 709318
rect 268502 709082 268586 709318
rect 268822 709082 268854 709318
rect 264514 707718 265134 707750
rect 264514 707482 264546 707718
rect 264782 707482 264866 707718
rect 265102 707482 265134 707718
rect 264514 707398 265134 707482
rect 264514 707162 264546 707398
rect 264782 707162 264866 707398
rect 265102 707162 265134 707398
rect 251954 693378 251986 693614
rect 252222 693378 252306 693614
rect 252542 693378 252574 693614
rect 251954 693294 252574 693378
rect 251954 693058 251986 693294
rect 252222 693058 252306 693294
rect 252542 693058 252574 693294
rect 251954 653614 252574 693058
rect 251954 653378 251986 653614
rect 252222 653378 252306 653614
rect 252542 653378 252574 653614
rect 251954 653294 252574 653378
rect 251954 653058 251986 653294
rect 252222 653058 252306 653294
rect 252542 653058 252574 653294
rect 251954 613614 252574 653058
rect 251954 613378 251986 613614
rect 252222 613378 252306 613614
rect 252542 613378 252574 613614
rect 251954 613294 252574 613378
rect 251954 613058 251986 613294
rect 252222 613058 252306 613294
rect 252542 613058 252574 613294
rect 251954 573614 252574 613058
rect 251954 573378 251986 573614
rect 252222 573378 252306 573614
rect 252542 573378 252574 573614
rect 251954 573294 252574 573378
rect 251954 573058 251986 573294
rect 252222 573058 252306 573294
rect 252542 573058 252574 573294
rect 251954 533614 252574 573058
rect 251954 533378 251986 533614
rect 252222 533378 252306 533614
rect 252542 533378 252574 533614
rect 251954 533294 252574 533378
rect 251954 533058 251986 533294
rect 252222 533058 252306 533294
rect 252542 533058 252574 533294
rect 251954 493614 252574 533058
rect 251954 493378 251986 493614
rect 252222 493378 252306 493614
rect 252542 493378 252574 493614
rect 251954 493294 252574 493378
rect 251954 493058 251986 493294
rect 252222 493058 252306 493294
rect 252542 493058 252574 493294
rect 251954 453614 252574 493058
rect 251954 453378 251986 453614
rect 252222 453378 252306 453614
rect 252542 453378 252574 453614
rect 251954 453294 252574 453378
rect 251954 453058 251986 453294
rect 252222 453058 252306 453294
rect 252542 453058 252574 453294
rect 251954 413614 252574 453058
rect 251954 413378 251986 413614
rect 252222 413378 252306 413614
rect 252542 413378 252574 413614
rect 251954 413294 252574 413378
rect 251954 413058 251986 413294
rect 252222 413058 252306 413294
rect 252542 413058 252574 413294
rect 251954 373614 252574 413058
rect 251954 373378 251986 373614
rect 252222 373378 252306 373614
rect 252542 373378 252574 373614
rect 251954 373294 252574 373378
rect 251954 373058 251986 373294
rect 252222 373058 252306 373294
rect 252542 373058 252574 373294
rect 251954 333614 252574 373058
rect 251954 333378 251986 333614
rect 252222 333378 252306 333614
rect 252542 333378 252574 333614
rect 251954 333294 252574 333378
rect 251954 333058 251986 333294
rect 252222 333058 252306 333294
rect 252542 333058 252574 333294
rect 251954 293614 252574 333058
rect 251954 293378 251986 293614
rect 252222 293378 252306 293614
rect 252542 293378 252574 293614
rect 251954 293294 252574 293378
rect 251954 293058 251986 293294
rect 252222 293058 252306 293294
rect 252542 293058 252574 293294
rect 251954 253614 252574 293058
rect 251954 253378 251986 253614
rect 252222 253378 252306 253614
rect 252542 253378 252574 253614
rect 251954 253294 252574 253378
rect 251954 253058 251986 253294
rect 252222 253058 252306 253294
rect 252542 253058 252574 253294
rect 251954 213614 252574 253058
rect 251954 213378 251986 213614
rect 252222 213378 252306 213614
rect 252542 213378 252574 213614
rect 251954 213294 252574 213378
rect 251954 213058 251986 213294
rect 252222 213058 252306 213294
rect 252542 213058 252574 213294
rect 251954 173614 252574 213058
rect 251954 173378 251986 173614
rect 252222 173378 252306 173614
rect 252542 173378 252574 173614
rect 251954 173294 252574 173378
rect 251954 173058 251986 173294
rect 252222 173058 252306 173294
rect 252542 173058 252574 173294
rect 251954 133614 252574 173058
rect 251954 133378 251986 133614
rect 252222 133378 252306 133614
rect 252542 133378 252574 133614
rect 251954 133294 252574 133378
rect 251954 133058 251986 133294
rect 252222 133058 252306 133294
rect 252542 133058 252574 133294
rect 251954 93614 252574 133058
rect 251954 93378 251986 93614
rect 252222 93378 252306 93614
rect 252542 93378 252574 93614
rect 251954 93294 252574 93378
rect 251954 93058 251986 93294
rect 252222 93058 252306 93294
rect 252542 93058 252574 93294
rect 251954 53614 252574 93058
rect 251954 53378 251986 53614
rect 252222 53378 252306 53614
rect 252542 53378 252574 53614
rect 251954 53294 252574 53378
rect 251954 53058 251986 53294
rect 252222 53058 252306 53294
rect 252542 53058 252574 53294
rect 251954 13614 252574 53058
rect 251954 13378 251986 13614
rect 252222 13378 252306 13614
rect 252542 13378 252574 13614
rect 251954 13294 252574 13378
rect 251954 13058 251986 13294
rect 252222 13058 252306 13294
rect 252542 13058 252574 13294
rect 231954 -7302 231986 -7066
rect 232222 -7302 232306 -7066
rect 232542 -7302 232574 -7066
rect 231954 -7386 232574 -7302
rect 231954 -7622 231986 -7386
rect 232222 -7622 232306 -7386
rect 232542 -7622 232574 -7386
rect 231954 -7654 232574 -7622
rect 251954 -6106 252574 13058
rect 260794 705798 261414 705830
rect 260794 705562 260826 705798
rect 261062 705562 261146 705798
rect 261382 705562 261414 705798
rect 260794 705478 261414 705562
rect 260794 705242 260826 705478
rect 261062 705242 261146 705478
rect 261382 705242 261414 705478
rect 260794 662454 261414 705242
rect 260794 662218 260826 662454
rect 261062 662218 261146 662454
rect 261382 662218 261414 662454
rect 260794 662134 261414 662218
rect 260794 661898 260826 662134
rect 261062 661898 261146 662134
rect 261382 661898 261414 662134
rect 260794 622454 261414 661898
rect 260794 622218 260826 622454
rect 261062 622218 261146 622454
rect 261382 622218 261414 622454
rect 260794 622134 261414 622218
rect 260794 621898 260826 622134
rect 261062 621898 261146 622134
rect 261382 621898 261414 622134
rect 260794 582454 261414 621898
rect 260794 582218 260826 582454
rect 261062 582218 261146 582454
rect 261382 582218 261414 582454
rect 260794 582134 261414 582218
rect 260794 581898 260826 582134
rect 261062 581898 261146 582134
rect 261382 581898 261414 582134
rect 260794 542454 261414 581898
rect 260794 542218 260826 542454
rect 261062 542218 261146 542454
rect 261382 542218 261414 542454
rect 260794 542134 261414 542218
rect 260794 541898 260826 542134
rect 261062 541898 261146 542134
rect 261382 541898 261414 542134
rect 260794 502454 261414 541898
rect 260794 502218 260826 502454
rect 261062 502218 261146 502454
rect 261382 502218 261414 502454
rect 260794 502134 261414 502218
rect 260794 501898 260826 502134
rect 261062 501898 261146 502134
rect 261382 501898 261414 502134
rect 260794 462454 261414 501898
rect 260794 462218 260826 462454
rect 261062 462218 261146 462454
rect 261382 462218 261414 462454
rect 260794 462134 261414 462218
rect 260794 461898 260826 462134
rect 261062 461898 261146 462134
rect 261382 461898 261414 462134
rect 260794 422454 261414 461898
rect 260794 422218 260826 422454
rect 261062 422218 261146 422454
rect 261382 422218 261414 422454
rect 260794 422134 261414 422218
rect 260794 421898 260826 422134
rect 261062 421898 261146 422134
rect 261382 421898 261414 422134
rect 260794 382454 261414 421898
rect 260794 382218 260826 382454
rect 261062 382218 261146 382454
rect 261382 382218 261414 382454
rect 260794 382134 261414 382218
rect 260794 381898 260826 382134
rect 261062 381898 261146 382134
rect 261382 381898 261414 382134
rect 260794 342454 261414 381898
rect 260794 342218 260826 342454
rect 261062 342218 261146 342454
rect 261382 342218 261414 342454
rect 260794 342134 261414 342218
rect 260794 341898 260826 342134
rect 261062 341898 261146 342134
rect 261382 341898 261414 342134
rect 260794 302454 261414 341898
rect 260794 302218 260826 302454
rect 261382 302218 261414 302454
rect 260794 302134 261414 302218
rect 260794 301898 260826 302134
rect 261382 301898 261414 302134
rect 260794 262454 261414 301898
rect 260794 262218 260826 262454
rect 261382 262218 261414 262454
rect 260794 262134 261414 262218
rect 260794 261898 260826 262134
rect 261382 261898 261414 262134
rect 260794 222454 261414 261898
rect 260794 222218 260826 222454
rect 261382 222218 261414 222454
rect 260794 222134 261414 222218
rect 260794 221898 260826 222134
rect 261382 221898 261414 222134
rect 260794 182454 261414 221898
rect 260794 182218 260826 182454
rect 261382 182218 261414 182454
rect 260794 182134 261414 182218
rect 260794 181898 260826 182134
rect 261382 181898 261414 182134
rect 260794 142454 261414 181898
rect 260794 142218 260826 142454
rect 261382 142218 261414 142454
rect 260794 142134 261414 142218
rect 260794 141898 260826 142134
rect 261382 141898 261414 142134
rect 260794 102454 261414 141898
rect 260794 102218 260826 102454
rect 261062 102218 261146 102454
rect 261382 102218 261414 102454
rect 260794 102134 261414 102218
rect 260794 101898 260826 102134
rect 261062 101898 261146 102134
rect 261382 101898 261414 102134
rect 260794 62454 261414 101898
rect 260794 62218 260826 62454
rect 261062 62218 261146 62454
rect 261382 62218 261414 62454
rect 260794 62134 261414 62218
rect 260794 61898 260826 62134
rect 261062 61898 261146 62134
rect 261382 61898 261414 62134
rect 260794 22454 261414 61898
rect 260794 22218 260826 22454
rect 261062 22218 261146 22454
rect 261382 22218 261414 22454
rect 260794 22134 261414 22218
rect 260794 21898 260826 22134
rect 261062 21898 261146 22134
rect 261382 21898 261414 22134
rect 260794 -1306 261414 21898
rect 260794 -1542 260826 -1306
rect 261062 -1542 261146 -1306
rect 261382 -1542 261414 -1306
rect 260794 -1626 261414 -1542
rect 260794 -1862 260826 -1626
rect 261062 -1862 261146 -1626
rect 261382 -1862 261414 -1626
rect 260794 -1894 261414 -1862
rect 264514 666174 265134 707162
rect 264514 665938 264546 666174
rect 264782 665938 264866 666174
rect 265102 665938 265134 666174
rect 264514 665854 265134 665938
rect 264514 665618 264546 665854
rect 264782 665618 264866 665854
rect 265102 665618 265134 665854
rect 264514 626174 265134 665618
rect 264514 625938 264546 626174
rect 264782 625938 264866 626174
rect 265102 625938 265134 626174
rect 264514 625854 265134 625938
rect 264514 625618 264546 625854
rect 264782 625618 264866 625854
rect 265102 625618 265134 625854
rect 264514 586174 265134 625618
rect 264514 585938 264546 586174
rect 264782 585938 264866 586174
rect 265102 585938 265134 586174
rect 264514 585854 265134 585938
rect 264514 585618 264546 585854
rect 264782 585618 264866 585854
rect 265102 585618 265134 585854
rect 264514 546174 265134 585618
rect 264514 545938 264546 546174
rect 264782 545938 264866 546174
rect 265102 545938 265134 546174
rect 264514 545854 265134 545938
rect 264514 545618 264546 545854
rect 264782 545618 264866 545854
rect 265102 545618 265134 545854
rect 264514 506174 265134 545618
rect 264514 505938 264546 506174
rect 264782 505938 264866 506174
rect 265102 505938 265134 506174
rect 264514 505854 265134 505938
rect 264514 505618 264546 505854
rect 264782 505618 264866 505854
rect 265102 505618 265134 505854
rect 264514 466174 265134 505618
rect 264514 465938 264546 466174
rect 264782 465938 264866 466174
rect 265102 465938 265134 466174
rect 264514 465854 265134 465938
rect 264514 465618 264546 465854
rect 264782 465618 264866 465854
rect 265102 465618 265134 465854
rect 264514 426174 265134 465618
rect 264514 425938 264546 426174
rect 264782 425938 264866 426174
rect 265102 425938 265134 426174
rect 264514 425854 265134 425938
rect 264514 425618 264546 425854
rect 264782 425618 264866 425854
rect 265102 425618 265134 425854
rect 264514 386174 265134 425618
rect 264514 385938 264546 386174
rect 264782 385938 264866 386174
rect 265102 385938 265134 386174
rect 264514 385854 265134 385938
rect 264514 385618 264546 385854
rect 264782 385618 264866 385854
rect 265102 385618 265134 385854
rect 264514 346174 265134 385618
rect 264514 345938 264546 346174
rect 264782 345938 264866 346174
rect 265102 345938 265134 346174
rect 264514 345854 265134 345938
rect 264514 345618 264546 345854
rect 264782 345618 264866 345854
rect 265102 345618 265134 345854
rect 264514 306174 265134 345618
rect 264514 305938 264546 306174
rect 264782 305938 264866 306174
rect 265102 305938 265134 306174
rect 264514 305854 265134 305938
rect 264514 305618 264546 305854
rect 264782 305618 264866 305854
rect 265102 305618 265134 305854
rect 264514 266174 265134 305618
rect 264514 265938 264546 266174
rect 264782 265938 264866 266174
rect 265102 265938 265134 266174
rect 264514 265854 265134 265938
rect 264514 265618 264546 265854
rect 264782 265618 264866 265854
rect 265102 265618 265134 265854
rect 264514 226174 265134 265618
rect 264514 225938 264546 226174
rect 264782 225938 264866 226174
rect 265102 225938 265134 226174
rect 264514 225854 265134 225938
rect 264514 225618 264546 225854
rect 264782 225618 264866 225854
rect 265102 225618 265134 225854
rect 264514 186174 265134 225618
rect 264514 185938 264546 186174
rect 264782 185938 264866 186174
rect 265102 185938 265134 186174
rect 264514 185854 265134 185938
rect 264514 185618 264546 185854
rect 264782 185618 264866 185854
rect 265102 185618 265134 185854
rect 264514 146174 265134 185618
rect 264514 145938 264546 146174
rect 264782 145938 264866 146174
rect 265102 145938 265134 146174
rect 264514 145854 265134 145938
rect 264514 145618 264546 145854
rect 264782 145618 264866 145854
rect 265102 145618 265134 145854
rect 264514 106174 265134 145618
rect 264514 105938 264546 106174
rect 264782 105938 264866 106174
rect 265102 105938 265134 106174
rect 264514 105854 265134 105938
rect 264514 105618 264546 105854
rect 264782 105618 264866 105854
rect 265102 105618 265134 105854
rect 264514 66174 265134 105618
rect 264514 65938 264546 66174
rect 264782 65938 264866 66174
rect 265102 65938 265134 66174
rect 264514 65854 265134 65938
rect 264514 65618 264546 65854
rect 264782 65618 264866 65854
rect 265102 65618 265134 65854
rect 264514 26174 265134 65618
rect 264514 25938 264546 26174
rect 264782 25938 264866 26174
rect 265102 25938 265134 26174
rect 264514 25854 265134 25938
rect 264514 25618 264546 25854
rect 264782 25618 264866 25854
rect 265102 25618 265134 25854
rect 264514 -3226 265134 25618
rect 264514 -3462 264546 -3226
rect 264782 -3462 264866 -3226
rect 265102 -3462 265134 -3226
rect 264514 -3546 265134 -3462
rect 264514 -3782 264546 -3546
rect 264782 -3782 264866 -3546
rect 265102 -3782 265134 -3546
rect 264514 -3814 265134 -3782
rect 268234 669894 268854 709082
rect 268234 669658 268266 669894
rect 268502 669658 268586 669894
rect 268822 669658 268854 669894
rect 268234 669574 268854 669658
rect 268234 669338 268266 669574
rect 268502 669338 268586 669574
rect 268822 669338 268854 669574
rect 268234 629894 268854 669338
rect 268234 629658 268266 629894
rect 268502 629658 268586 629894
rect 268822 629658 268854 629894
rect 268234 629574 268854 629658
rect 268234 629338 268266 629574
rect 268502 629338 268586 629574
rect 268822 629338 268854 629574
rect 268234 589894 268854 629338
rect 268234 589658 268266 589894
rect 268502 589658 268586 589894
rect 268822 589658 268854 589894
rect 268234 589574 268854 589658
rect 268234 589338 268266 589574
rect 268502 589338 268586 589574
rect 268822 589338 268854 589574
rect 268234 549894 268854 589338
rect 268234 549658 268266 549894
rect 268502 549658 268586 549894
rect 268822 549658 268854 549894
rect 268234 549574 268854 549658
rect 268234 549338 268266 549574
rect 268502 549338 268586 549574
rect 268822 549338 268854 549574
rect 268234 509894 268854 549338
rect 268234 509658 268266 509894
rect 268502 509658 268586 509894
rect 268822 509658 268854 509894
rect 268234 509574 268854 509658
rect 268234 509338 268266 509574
rect 268502 509338 268586 509574
rect 268822 509338 268854 509574
rect 268234 469894 268854 509338
rect 268234 469658 268266 469894
rect 268502 469658 268586 469894
rect 268822 469658 268854 469894
rect 268234 469574 268854 469658
rect 268234 469338 268266 469574
rect 268502 469338 268586 469574
rect 268822 469338 268854 469574
rect 268234 429894 268854 469338
rect 268234 429658 268266 429894
rect 268502 429658 268586 429894
rect 268822 429658 268854 429894
rect 268234 429574 268854 429658
rect 268234 429338 268266 429574
rect 268502 429338 268586 429574
rect 268822 429338 268854 429574
rect 268234 389894 268854 429338
rect 268234 389658 268266 389894
rect 268502 389658 268586 389894
rect 268822 389658 268854 389894
rect 268234 389574 268854 389658
rect 268234 389338 268266 389574
rect 268502 389338 268586 389574
rect 268822 389338 268854 389574
rect 268234 349894 268854 389338
rect 268234 349658 268266 349894
rect 268502 349658 268586 349894
rect 268822 349658 268854 349894
rect 268234 349574 268854 349658
rect 268234 349338 268266 349574
rect 268502 349338 268586 349574
rect 268822 349338 268854 349574
rect 268234 309894 268854 349338
rect 268234 309658 268266 309894
rect 268502 309658 268586 309894
rect 268822 309658 268854 309894
rect 268234 309574 268854 309658
rect 268234 309338 268266 309574
rect 268502 309338 268586 309574
rect 268822 309338 268854 309574
rect 268234 269894 268854 309338
rect 268234 269658 268266 269894
rect 268502 269658 268586 269894
rect 268822 269658 268854 269894
rect 268234 269574 268854 269658
rect 268234 269338 268266 269574
rect 268502 269338 268586 269574
rect 268822 269338 268854 269574
rect 268234 229894 268854 269338
rect 268234 229658 268266 229894
rect 268502 229658 268586 229894
rect 268822 229658 268854 229894
rect 268234 229574 268854 229658
rect 268234 229338 268266 229574
rect 268502 229338 268586 229574
rect 268822 229338 268854 229574
rect 268234 189894 268854 229338
rect 268234 189658 268266 189894
rect 268502 189658 268586 189894
rect 268822 189658 268854 189894
rect 268234 189574 268854 189658
rect 268234 189338 268266 189574
rect 268502 189338 268586 189574
rect 268822 189338 268854 189574
rect 268234 149894 268854 189338
rect 268234 149658 268266 149894
rect 268502 149658 268586 149894
rect 268822 149658 268854 149894
rect 268234 149574 268854 149658
rect 268234 149338 268266 149574
rect 268502 149338 268586 149574
rect 268822 149338 268854 149574
rect 268234 109894 268854 149338
rect 268234 109658 268266 109894
rect 268502 109658 268586 109894
rect 268822 109658 268854 109894
rect 268234 109574 268854 109658
rect 268234 109338 268266 109574
rect 268502 109338 268586 109574
rect 268822 109338 268854 109574
rect 268234 69894 268854 109338
rect 268234 69658 268266 69894
rect 268502 69658 268586 69894
rect 268822 69658 268854 69894
rect 268234 69574 268854 69658
rect 268234 69338 268266 69574
rect 268502 69338 268586 69574
rect 268822 69338 268854 69574
rect 268234 29894 268854 69338
rect 268234 29658 268266 29894
rect 268502 29658 268586 29894
rect 268822 29658 268854 29894
rect 268234 29574 268854 29658
rect 268234 29338 268266 29574
rect 268502 29338 268586 29574
rect 268822 29338 268854 29574
rect 268234 -5146 268854 29338
rect 268234 -5382 268266 -5146
rect 268502 -5382 268586 -5146
rect 268822 -5382 268854 -5146
rect 268234 -5466 268854 -5382
rect 268234 -5702 268266 -5466
rect 268502 -5702 268586 -5466
rect 268822 -5702 268854 -5466
rect 268234 -5734 268854 -5702
rect 271954 673614 272574 711002
rect 291954 710598 292574 711590
rect 291954 710362 291986 710598
rect 292222 710362 292306 710598
rect 292542 710362 292574 710598
rect 291954 710278 292574 710362
rect 291954 710042 291986 710278
rect 292222 710042 292306 710278
rect 292542 710042 292574 710278
rect 288234 708678 288854 709670
rect 288234 708442 288266 708678
rect 288502 708442 288586 708678
rect 288822 708442 288854 708678
rect 288234 708358 288854 708442
rect 288234 708122 288266 708358
rect 288502 708122 288586 708358
rect 288822 708122 288854 708358
rect 284514 706758 285134 707750
rect 284514 706522 284546 706758
rect 284782 706522 284866 706758
rect 285102 706522 285134 706758
rect 284514 706438 285134 706522
rect 284514 706202 284546 706438
rect 284782 706202 284866 706438
rect 285102 706202 285134 706438
rect 271954 673378 271986 673614
rect 272222 673378 272306 673614
rect 272542 673378 272574 673614
rect 271954 673294 272574 673378
rect 271954 673058 271986 673294
rect 272222 673058 272306 673294
rect 272542 673058 272574 673294
rect 271954 633614 272574 673058
rect 271954 633378 271986 633614
rect 272222 633378 272306 633614
rect 272542 633378 272574 633614
rect 271954 633294 272574 633378
rect 271954 633058 271986 633294
rect 272222 633058 272306 633294
rect 272542 633058 272574 633294
rect 271954 593614 272574 633058
rect 271954 593378 271986 593614
rect 272222 593378 272306 593614
rect 272542 593378 272574 593614
rect 271954 593294 272574 593378
rect 271954 593058 271986 593294
rect 272222 593058 272306 593294
rect 272542 593058 272574 593294
rect 271954 553614 272574 593058
rect 271954 553378 271986 553614
rect 272222 553378 272306 553614
rect 272542 553378 272574 553614
rect 271954 553294 272574 553378
rect 271954 553058 271986 553294
rect 272222 553058 272306 553294
rect 272542 553058 272574 553294
rect 271954 513614 272574 553058
rect 271954 513378 271986 513614
rect 272222 513378 272306 513614
rect 272542 513378 272574 513614
rect 271954 513294 272574 513378
rect 271954 513058 271986 513294
rect 272222 513058 272306 513294
rect 272542 513058 272574 513294
rect 271954 473614 272574 513058
rect 271954 473378 271986 473614
rect 272222 473378 272306 473614
rect 272542 473378 272574 473614
rect 271954 473294 272574 473378
rect 271954 473058 271986 473294
rect 272222 473058 272306 473294
rect 272542 473058 272574 473294
rect 271954 433614 272574 473058
rect 271954 433378 271986 433614
rect 272222 433378 272306 433614
rect 272542 433378 272574 433614
rect 271954 433294 272574 433378
rect 271954 433058 271986 433294
rect 272222 433058 272306 433294
rect 272542 433058 272574 433294
rect 271954 393614 272574 433058
rect 271954 393378 271986 393614
rect 272222 393378 272306 393614
rect 272542 393378 272574 393614
rect 271954 393294 272574 393378
rect 271954 393058 271986 393294
rect 272222 393058 272306 393294
rect 272542 393058 272574 393294
rect 271954 353614 272574 393058
rect 271954 353378 271986 353614
rect 272222 353378 272306 353614
rect 272542 353378 272574 353614
rect 271954 353294 272574 353378
rect 271954 353058 271986 353294
rect 272222 353058 272306 353294
rect 272542 353058 272574 353294
rect 271954 313614 272574 353058
rect 280794 704838 281414 705830
rect 280794 704602 280826 704838
rect 281062 704602 281146 704838
rect 281382 704602 281414 704838
rect 280794 704518 281414 704602
rect 280794 704282 280826 704518
rect 281062 704282 281146 704518
rect 281382 704282 281414 704518
rect 280794 682454 281414 704282
rect 280794 682218 280826 682454
rect 281062 682218 281146 682454
rect 281382 682218 281414 682454
rect 280794 682134 281414 682218
rect 280794 681898 280826 682134
rect 281062 681898 281146 682134
rect 281382 681898 281414 682134
rect 280794 642454 281414 681898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 602454 281414 641898
rect 280794 602218 280826 602454
rect 281062 602218 281146 602454
rect 281382 602218 281414 602454
rect 280794 602134 281414 602218
rect 280794 601898 280826 602134
rect 281062 601898 281146 602134
rect 281382 601898 281414 602134
rect 280794 562454 281414 601898
rect 280794 562218 280826 562454
rect 281062 562218 281146 562454
rect 281382 562218 281414 562454
rect 280794 562134 281414 562218
rect 280794 561898 280826 562134
rect 281062 561898 281146 562134
rect 281382 561898 281414 562134
rect 280794 522454 281414 561898
rect 280794 522218 280826 522454
rect 281062 522218 281146 522454
rect 281382 522218 281414 522454
rect 280794 522134 281414 522218
rect 280794 521898 280826 522134
rect 281062 521898 281146 522134
rect 281382 521898 281414 522134
rect 280794 482454 281414 521898
rect 280794 482218 280826 482454
rect 281062 482218 281146 482454
rect 281382 482218 281414 482454
rect 280794 482134 281414 482218
rect 280794 481898 280826 482134
rect 281062 481898 281146 482134
rect 281382 481898 281414 482134
rect 280794 442454 281414 481898
rect 280794 442218 280826 442454
rect 281062 442218 281146 442454
rect 281382 442218 281414 442454
rect 280794 442134 281414 442218
rect 280794 441898 280826 442134
rect 281062 441898 281146 442134
rect 281382 441898 281414 442134
rect 280794 402454 281414 441898
rect 280794 402218 280826 402454
rect 281062 402218 281146 402454
rect 281382 402218 281414 402454
rect 280794 402134 281414 402218
rect 280794 401898 280826 402134
rect 281062 401898 281146 402134
rect 281382 401898 281414 402134
rect 280794 362454 281414 401898
rect 280794 362218 280826 362454
rect 281062 362218 281146 362454
rect 281382 362218 281414 362454
rect 280794 362134 281414 362218
rect 280794 361898 280826 362134
rect 281062 361898 281146 362134
rect 281382 361898 281414 362134
rect 280794 322454 281414 361898
rect 280794 322218 280826 322454
rect 281062 322218 281146 322454
rect 281382 322218 281414 322454
rect 280794 322134 281414 322218
rect 280794 321898 280826 322134
rect 281062 321898 281146 322134
rect 281382 321898 281414 322134
rect 273299 319428 273365 319429
rect 273299 319364 273300 319428
rect 273364 319364 273365 319428
rect 273299 319363 273365 319364
rect 271954 313378 271986 313614
rect 272222 313378 272306 313614
rect 272542 313378 272574 313614
rect 271954 313294 272574 313378
rect 271954 313058 271986 313294
rect 272222 313058 272306 313294
rect 272542 313058 272574 313294
rect 271954 273614 272574 313058
rect 271954 273378 271986 273614
rect 272222 273378 272306 273614
rect 272542 273378 272574 273614
rect 271954 273294 272574 273378
rect 271954 273058 271986 273294
rect 272222 273058 272306 273294
rect 272542 273058 272574 273294
rect 271954 233614 272574 273058
rect 271954 233378 271986 233614
rect 272222 233378 272306 233614
rect 272542 233378 272574 233614
rect 271954 233294 272574 233378
rect 271954 233058 271986 233294
rect 272222 233058 272306 233294
rect 272542 233058 272574 233294
rect 271954 193614 272574 233058
rect 271954 193378 271986 193614
rect 272222 193378 272306 193614
rect 272542 193378 272574 193614
rect 271954 193294 272574 193378
rect 271954 193058 271986 193294
rect 272222 193058 272306 193294
rect 272542 193058 272574 193294
rect 271954 153614 272574 193058
rect 271954 153378 271986 153614
rect 272222 153378 272306 153614
rect 272542 153378 272574 153614
rect 271954 153294 272574 153378
rect 271954 153058 271986 153294
rect 272222 153058 272306 153294
rect 272542 153058 272574 153294
rect 271954 113614 272574 153058
rect 271954 113378 271986 113614
rect 272222 113378 272306 113614
rect 272542 113378 272574 113614
rect 271954 113294 272574 113378
rect 271954 113058 271986 113294
rect 272222 113058 272306 113294
rect 272542 113058 272574 113294
rect 271954 73614 272574 113058
rect 271954 73378 271986 73614
rect 272222 73378 272306 73614
rect 272542 73378 272574 73614
rect 271954 73294 272574 73378
rect 271954 73058 271986 73294
rect 272222 73058 272306 73294
rect 272542 73058 272574 73294
rect 271954 33614 272574 73058
rect 271954 33378 271986 33614
rect 272222 33378 272306 33614
rect 272542 33378 272574 33614
rect 271954 33294 272574 33378
rect 271954 33058 271986 33294
rect 272222 33058 272306 33294
rect 272542 33058 272574 33294
rect 251954 -6342 251986 -6106
rect 252222 -6342 252306 -6106
rect 252542 -6342 252574 -6106
rect 251954 -6426 252574 -6342
rect 251954 -6662 251986 -6426
rect 252222 -6662 252306 -6426
rect 252542 -6662 252574 -6426
rect 251954 -7654 252574 -6662
rect 271954 -7066 272574 33058
rect 273302 3773 273362 319363
rect 280794 282454 281414 321898
rect 284514 686174 285134 706202
rect 284514 685938 284546 686174
rect 284782 685938 284866 686174
rect 285102 685938 285134 686174
rect 284514 685854 285134 685938
rect 284514 685618 284546 685854
rect 284782 685618 284866 685854
rect 285102 685618 285134 685854
rect 284514 646174 285134 685618
rect 284514 645938 284546 646174
rect 284782 645938 284866 646174
rect 285102 645938 285134 646174
rect 284514 645854 285134 645938
rect 284514 645618 284546 645854
rect 284782 645618 284866 645854
rect 285102 645618 285134 645854
rect 284514 606174 285134 645618
rect 284514 605938 284546 606174
rect 284782 605938 284866 606174
rect 285102 605938 285134 606174
rect 284514 605854 285134 605938
rect 284514 605618 284546 605854
rect 284782 605618 284866 605854
rect 285102 605618 285134 605854
rect 284514 566174 285134 605618
rect 284514 565938 284546 566174
rect 284782 565938 284866 566174
rect 285102 565938 285134 566174
rect 284514 565854 285134 565938
rect 284514 565618 284546 565854
rect 284782 565618 284866 565854
rect 285102 565618 285134 565854
rect 284514 526174 285134 565618
rect 284514 525938 284546 526174
rect 284782 525938 284866 526174
rect 285102 525938 285134 526174
rect 284514 525854 285134 525938
rect 284514 525618 284546 525854
rect 284782 525618 284866 525854
rect 285102 525618 285134 525854
rect 284514 486174 285134 525618
rect 284514 485938 284546 486174
rect 284782 485938 284866 486174
rect 285102 485938 285134 486174
rect 284514 485854 285134 485938
rect 284514 485618 284546 485854
rect 284782 485618 284866 485854
rect 285102 485618 285134 485854
rect 284514 446174 285134 485618
rect 284514 445938 284546 446174
rect 284782 445938 284866 446174
rect 285102 445938 285134 446174
rect 284514 445854 285134 445938
rect 284514 445618 284546 445854
rect 284782 445618 284866 445854
rect 285102 445618 285134 445854
rect 284514 406174 285134 445618
rect 284514 405938 284546 406174
rect 284782 405938 284866 406174
rect 285102 405938 285134 406174
rect 284514 405854 285134 405938
rect 284514 405618 284546 405854
rect 284782 405618 284866 405854
rect 285102 405618 285134 405854
rect 284514 366174 285134 405618
rect 284514 365938 284546 366174
rect 284782 365938 284866 366174
rect 285102 365938 285134 366174
rect 284514 365854 285134 365938
rect 284514 365618 284546 365854
rect 284782 365618 284866 365854
rect 285102 365618 285134 365854
rect 284514 326174 285134 365618
rect 284514 325938 284546 326174
rect 284782 325938 284866 326174
rect 285102 325938 285134 326174
rect 284514 325854 285134 325938
rect 284514 325618 284546 325854
rect 284782 325618 284866 325854
rect 285102 325618 285134 325854
rect 282867 319428 282933 319429
rect 282867 319364 282868 319428
rect 282932 319364 282933 319428
rect 282867 319363 282933 319364
rect 280794 282218 280826 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281382 281898 281414 282134
rect 280794 242454 281414 281898
rect 280794 242218 280826 242454
rect 281382 242218 281414 242454
rect 280794 242134 281414 242218
rect 280794 241898 280826 242134
rect 281382 241898 281414 242134
rect 280794 202454 281414 241898
rect 280794 202218 280826 202454
rect 281382 202218 281414 202454
rect 280794 202134 281414 202218
rect 280794 201898 280826 202134
rect 281382 201898 281414 202134
rect 280794 162454 281414 201898
rect 280794 162218 280826 162454
rect 281382 162218 281414 162454
rect 280794 162134 281414 162218
rect 280794 161898 280826 162134
rect 281382 161898 281414 162134
rect 280794 122454 281414 161898
rect 280794 122218 280826 122454
rect 281062 122218 281146 122454
rect 281382 122218 281414 122454
rect 280794 122134 281414 122218
rect 280794 121898 280826 122134
rect 281062 121898 281146 122134
rect 281382 121898 281414 122134
rect 280794 82454 281414 121898
rect 280794 82218 280826 82454
rect 281062 82218 281146 82454
rect 281382 82218 281414 82454
rect 280794 82134 281414 82218
rect 280794 81898 280826 82134
rect 281062 81898 281146 82134
rect 281382 81898 281414 82134
rect 280794 42454 281414 81898
rect 280794 42218 280826 42454
rect 281062 42218 281146 42454
rect 281382 42218 281414 42454
rect 280794 42134 281414 42218
rect 280794 41898 280826 42134
rect 281062 41898 281146 42134
rect 281382 41898 281414 42134
rect 273299 3772 273365 3773
rect 273299 3708 273300 3772
rect 273364 3708 273365 3772
rect 273299 3707 273365 3708
rect 280794 2454 281414 41898
rect 282870 3501 282930 319363
rect 284514 286174 285134 325618
rect 284514 285938 284546 286174
rect 284782 285938 284866 286174
rect 285102 285938 285134 286174
rect 284514 285854 285134 285938
rect 284514 285618 284546 285854
rect 284782 285618 284866 285854
rect 285102 285618 285134 285854
rect 284514 246174 285134 285618
rect 284514 245938 284546 246174
rect 284782 245938 284866 246174
rect 285102 245938 285134 246174
rect 284514 245854 285134 245938
rect 284514 245618 284546 245854
rect 284782 245618 284866 245854
rect 285102 245618 285134 245854
rect 284514 206174 285134 245618
rect 284514 205938 284546 206174
rect 284782 205938 284866 206174
rect 285102 205938 285134 206174
rect 284514 205854 285134 205938
rect 284514 205618 284546 205854
rect 284782 205618 284866 205854
rect 285102 205618 285134 205854
rect 284514 166174 285134 205618
rect 284514 165938 284546 166174
rect 284782 165938 284866 166174
rect 285102 165938 285134 166174
rect 284514 165854 285134 165938
rect 284514 165618 284546 165854
rect 284782 165618 284866 165854
rect 285102 165618 285134 165854
rect 284514 126174 285134 165618
rect 284514 125938 284546 126174
rect 284782 125938 284866 126174
rect 285102 125938 285134 126174
rect 284514 125854 285134 125938
rect 284514 125618 284546 125854
rect 284782 125618 284866 125854
rect 285102 125618 285134 125854
rect 284514 86174 285134 125618
rect 284514 85938 284546 86174
rect 284782 85938 284866 86174
rect 285102 85938 285134 86174
rect 284514 85854 285134 85938
rect 284514 85618 284546 85854
rect 284782 85618 284866 85854
rect 285102 85618 285134 85854
rect 284514 46174 285134 85618
rect 284514 45938 284546 46174
rect 284782 45938 284866 46174
rect 285102 45938 285134 46174
rect 284514 45854 285134 45938
rect 284514 45618 284546 45854
rect 284782 45618 284866 45854
rect 285102 45618 285134 45854
rect 284514 6174 285134 45618
rect 284514 5938 284546 6174
rect 284782 5938 284866 6174
rect 285102 5938 285134 6174
rect 284514 5854 285134 5938
rect 284514 5618 284546 5854
rect 284782 5618 284866 5854
rect 285102 5618 285134 5854
rect 282867 3500 282933 3501
rect 282867 3436 282868 3500
rect 282932 3436 282933 3500
rect 282867 3435 282933 3436
rect 280794 2218 280826 2454
rect 281062 2218 281146 2454
rect 281382 2218 281414 2454
rect 280794 2134 281414 2218
rect 280794 1898 280826 2134
rect 281062 1898 281146 2134
rect 281382 1898 281414 2134
rect 280794 -346 281414 1898
rect 280794 -582 280826 -346
rect 281062 -582 281146 -346
rect 281382 -582 281414 -346
rect 280794 -666 281414 -582
rect 280794 -902 280826 -666
rect 281062 -902 281146 -666
rect 281382 -902 281414 -666
rect 280794 -1894 281414 -902
rect 284514 -2266 285134 5618
rect 284514 -2502 284546 -2266
rect 284782 -2502 284866 -2266
rect 285102 -2502 285134 -2266
rect 284514 -2586 285134 -2502
rect 284514 -2822 284546 -2586
rect 284782 -2822 284866 -2586
rect 285102 -2822 285134 -2586
rect 284514 -3814 285134 -2822
rect 288234 689894 288854 708122
rect 288234 689658 288266 689894
rect 288502 689658 288586 689894
rect 288822 689658 288854 689894
rect 288234 689574 288854 689658
rect 288234 689338 288266 689574
rect 288502 689338 288586 689574
rect 288822 689338 288854 689574
rect 288234 649894 288854 689338
rect 288234 649658 288266 649894
rect 288502 649658 288586 649894
rect 288822 649658 288854 649894
rect 288234 649574 288854 649658
rect 288234 649338 288266 649574
rect 288502 649338 288586 649574
rect 288822 649338 288854 649574
rect 288234 609894 288854 649338
rect 288234 609658 288266 609894
rect 288502 609658 288586 609894
rect 288822 609658 288854 609894
rect 288234 609574 288854 609658
rect 288234 609338 288266 609574
rect 288502 609338 288586 609574
rect 288822 609338 288854 609574
rect 288234 569894 288854 609338
rect 288234 569658 288266 569894
rect 288502 569658 288586 569894
rect 288822 569658 288854 569894
rect 288234 569574 288854 569658
rect 288234 569338 288266 569574
rect 288502 569338 288586 569574
rect 288822 569338 288854 569574
rect 288234 529894 288854 569338
rect 288234 529658 288266 529894
rect 288502 529658 288586 529894
rect 288822 529658 288854 529894
rect 288234 529574 288854 529658
rect 288234 529338 288266 529574
rect 288502 529338 288586 529574
rect 288822 529338 288854 529574
rect 288234 489894 288854 529338
rect 288234 489658 288266 489894
rect 288502 489658 288586 489894
rect 288822 489658 288854 489894
rect 288234 489574 288854 489658
rect 288234 489338 288266 489574
rect 288502 489338 288586 489574
rect 288822 489338 288854 489574
rect 288234 449894 288854 489338
rect 288234 449658 288266 449894
rect 288502 449658 288586 449894
rect 288822 449658 288854 449894
rect 288234 449574 288854 449658
rect 288234 449338 288266 449574
rect 288502 449338 288586 449574
rect 288822 449338 288854 449574
rect 288234 409894 288854 449338
rect 288234 409658 288266 409894
rect 288502 409658 288586 409894
rect 288822 409658 288854 409894
rect 288234 409574 288854 409658
rect 288234 409338 288266 409574
rect 288502 409338 288586 409574
rect 288822 409338 288854 409574
rect 288234 369894 288854 409338
rect 288234 369658 288266 369894
rect 288502 369658 288586 369894
rect 288822 369658 288854 369894
rect 288234 369574 288854 369658
rect 288234 369338 288266 369574
rect 288502 369338 288586 369574
rect 288822 369338 288854 369574
rect 288234 329894 288854 369338
rect 288234 329658 288266 329894
rect 288502 329658 288586 329894
rect 288822 329658 288854 329894
rect 288234 329574 288854 329658
rect 288234 329338 288266 329574
rect 288502 329338 288586 329574
rect 288822 329338 288854 329574
rect 288234 289894 288854 329338
rect 288234 289658 288266 289894
rect 288502 289658 288586 289894
rect 288822 289658 288854 289894
rect 288234 289574 288854 289658
rect 288234 289338 288266 289574
rect 288502 289338 288586 289574
rect 288822 289338 288854 289574
rect 288234 249894 288854 289338
rect 288234 249658 288266 249894
rect 288502 249658 288586 249894
rect 288822 249658 288854 249894
rect 288234 249574 288854 249658
rect 288234 249338 288266 249574
rect 288502 249338 288586 249574
rect 288822 249338 288854 249574
rect 288234 209894 288854 249338
rect 288234 209658 288266 209894
rect 288502 209658 288586 209894
rect 288822 209658 288854 209894
rect 288234 209574 288854 209658
rect 288234 209338 288266 209574
rect 288502 209338 288586 209574
rect 288822 209338 288854 209574
rect 288234 169894 288854 209338
rect 288234 169658 288266 169894
rect 288502 169658 288586 169894
rect 288822 169658 288854 169894
rect 288234 169574 288854 169658
rect 288234 169338 288266 169574
rect 288502 169338 288586 169574
rect 288822 169338 288854 169574
rect 288234 129894 288854 169338
rect 288234 129658 288266 129894
rect 288502 129658 288586 129894
rect 288822 129658 288854 129894
rect 288234 129574 288854 129658
rect 288234 129338 288266 129574
rect 288502 129338 288586 129574
rect 288822 129338 288854 129574
rect 288234 89894 288854 129338
rect 288234 89658 288266 89894
rect 288502 89658 288586 89894
rect 288822 89658 288854 89894
rect 288234 89574 288854 89658
rect 288234 89338 288266 89574
rect 288502 89338 288586 89574
rect 288822 89338 288854 89574
rect 288234 49894 288854 89338
rect 288234 49658 288266 49894
rect 288502 49658 288586 49894
rect 288822 49658 288854 49894
rect 288234 49574 288854 49658
rect 288234 49338 288266 49574
rect 288502 49338 288586 49574
rect 288822 49338 288854 49574
rect 288234 9894 288854 49338
rect 288234 9658 288266 9894
rect 288502 9658 288586 9894
rect 288822 9658 288854 9894
rect 288234 9574 288854 9658
rect 288234 9338 288266 9574
rect 288502 9338 288586 9574
rect 288822 9338 288854 9574
rect 288234 -4186 288854 9338
rect 288234 -4422 288266 -4186
rect 288502 -4422 288586 -4186
rect 288822 -4422 288854 -4186
rect 288234 -4506 288854 -4422
rect 288234 -4742 288266 -4506
rect 288502 -4742 288586 -4506
rect 288822 -4742 288854 -4506
rect 288234 -5734 288854 -4742
rect 291954 693614 292574 710042
rect 311954 711558 312574 711590
rect 311954 711322 311986 711558
rect 312222 711322 312306 711558
rect 312542 711322 312574 711558
rect 311954 711238 312574 711322
rect 311954 711002 311986 711238
rect 312222 711002 312306 711238
rect 312542 711002 312574 711238
rect 308234 709638 308854 709670
rect 308234 709402 308266 709638
rect 308502 709402 308586 709638
rect 308822 709402 308854 709638
rect 308234 709318 308854 709402
rect 308234 709082 308266 709318
rect 308502 709082 308586 709318
rect 308822 709082 308854 709318
rect 304514 707718 305134 707750
rect 304514 707482 304546 707718
rect 304782 707482 304866 707718
rect 305102 707482 305134 707718
rect 304514 707398 305134 707482
rect 304514 707162 304546 707398
rect 304782 707162 304866 707398
rect 305102 707162 305134 707398
rect 291954 693378 291986 693614
rect 292222 693378 292306 693614
rect 292542 693378 292574 693614
rect 291954 693294 292574 693378
rect 291954 693058 291986 693294
rect 292222 693058 292306 693294
rect 292542 693058 292574 693294
rect 291954 653614 292574 693058
rect 291954 653378 291986 653614
rect 292222 653378 292306 653614
rect 292542 653378 292574 653614
rect 291954 653294 292574 653378
rect 291954 653058 291986 653294
rect 292222 653058 292306 653294
rect 292542 653058 292574 653294
rect 291954 613614 292574 653058
rect 291954 613378 291986 613614
rect 292222 613378 292306 613614
rect 292542 613378 292574 613614
rect 291954 613294 292574 613378
rect 291954 613058 291986 613294
rect 292222 613058 292306 613294
rect 292542 613058 292574 613294
rect 291954 573614 292574 613058
rect 291954 573378 291986 573614
rect 292222 573378 292306 573614
rect 292542 573378 292574 573614
rect 291954 573294 292574 573378
rect 291954 573058 291986 573294
rect 292222 573058 292306 573294
rect 292542 573058 292574 573294
rect 291954 533614 292574 573058
rect 291954 533378 291986 533614
rect 292222 533378 292306 533614
rect 292542 533378 292574 533614
rect 291954 533294 292574 533378
rect 291954 533058 291986 533294
rect 292222 533058 292306 533294
rect 292542 533058 292574 533294
rect 291954 493614 292574 533058
rect 291954 493378 291986 493614
rect 292222 493378 292306 493614
rect 292542 493378 292574 493614
rect 291954 493294 292574 493378
rect 291954 493058 291986 493294
rect 292222 493058 292306 493294
rect 292542 493058 292574 493294
rect 291954 453614 292574 493058
rect 291954 453378 291986 453614
rect 292222 453378 292306 453614
rect 292542 453378 292574 453614
rect 291954 453294 292574 453378
rect 291954 453058 291986 453294
rect 292222 453058 292306 453294
rect 292542 453058 292574 453294
rect 291954 413614 292574 453058
rect 291954 413378 291986 413614
rect 292222 413378 292306 413614
rect 292542 413378 292574 413614
rect 291954 413294 292574 413378
rect 291954 413058 291986 413294
rect 292222 413058 292306 413294
rect 292542 413058 292574 413294
rect 291954 373614 292574 413058
rect 291954 373378 291986 373614
rect 292222 373378 292306 373614
rect 292542 373378 292574 373614
rect 291954 373294 292574 373378
rect 291954 373058 291986 373294
rect 292222 373058 292306 373294
rect 292542 373058 292574 373294
rect 291954 333614 292574 373058
rect 291954 333378 291986 333614
rect 292222 333378 292306 333614
rect 292542 333378 292574 333614
rect 291954 333294 292574 333378
rect 291954 333058 291986 333294
rect 292222 333058 292306 333294
rect 292542 333058 292574 333294
rect 291954 293614 292574 333058
rect 300794 705798 301414 705830
rect 300794 705562 300826 705798
rect 301062 705562 301146 705798
rect 301382 705562 301414 705798
rect 300794 705478 301414 705562
rect 300794 705242 300826 705478
rect 301062 705242 301146 705478
rect 301382 705242 301414 705478
rect 300794 662454 301414 705242
rect 300794 662218 300826 662454
rect 301062 662218 301146 662454
rect 301382 662218 301414 662454
rect 300794 662134 301414 662218
rect 300794 661898 300826 662134
rect 301062 661898 301146 662134
rect 301382 661898 301414 662134
rect 300794 622454 301414 661898
rect 300794 622218 300826 622454
rect 301062 622218 301146 622454
rect 301382 622218 301414 622454
rect 300794 622134 301414 622218
rect 300794 621898 300826 622134
rect 301062 621898 301146 622134
rect 301382 621898 301414 622134
rect 300794 582454 301414 621898
rect 300794 582218 300826 582454
rect 301062 582218 301146 582454
rect 301382 582218 301414 582454
rect 300794 582134 301414 582218
rect 300794 581898 300826 582134
rect 301062 581898 301146 582134
rect 301382 581898 301414 582134
rect 300794 542454 301414 581898
rect 300794 542218 300826 542454
rect 301062 542218 301146 542454
rect 301382 542218 301414 542454
rect 300794 542134 301414 542218
rect 300794 541898 300826 542134
rect 301062 541898 301146 542134
rect 301382 541898 301414 542134
rect 300794 502454 301414 541898
rect 300794 502218 300826 502454
rect 301062 502218 301146 502454
rect 301382 502218 301414 502454
rect 300794 502134 301414 502218
rect 300794 501898 300826 502134
rect 301062 501898 301146 502134
rect 301382 501898 301414 502134
rect 300794 462454 301414 501898
rect 300794 462218 300826 462454
rect 301062 462218 301146 462454
rect 301382 462218 301414 462454
rect 300794 462134 301414 462218
rect 300794 461898 300826 462134
rect 301062 461898 301146 462134
rect 301382 461898 301414 462134
rect 300794 422454 301414 461898
rect 300794 422218 300826 422454
rect 301062 422218 301146 422454
rect 301382 422218 301414 422454
rect 300794 422134 301414 422218
rect 300794 421898 300826 422134
rect 301062 421898 301146 422134
rect 301382 421898 301414 422134
rect 300794 382454 301414 421898
rect 300794 382218 300826 382454
rect 301062 382218 301146 382454
rect 301382 382218 301414 382454
rect 300794 382134 301414 382218
rect 300794 381898 300826 382134
rect 301062 381898 301146 382134
rect 301382 381898 301414 382134
rect 300794 342454 301414 381898
rect 300794 342218 300826 342454
rect 301062 342218 301146 342454
rect 301382 342218 301414 342454
rect 300794 342134 301414 342218
rect 300794 341898 300826 342134
rect 301062 341898 301146 342134
rect 301382 341898 301414 342134
rect 293907 319428 293973 319429
rect 293907 319364 293908 319428
rect 293972 319364 293973 319428
rect 293907 319363 293973 319364
rect 291954 293378 291986 293614
rect 292222 293378 292306 293614
rect 292542 293378 292574 293614
rect 291954 293294 292574 293378
rect 291954 293058 291986 293294
rect 292222 293058 292306 293294
rect 292542 293058 292574 293294
rect 291954 253614 292574 293058
rect 291954 253378 291986 253614
rect 292222 253378 292306 253614
rect 292542 253378 292574 253614
rect 291954 253294 292574 253378
rect 291954 253058 291986 253294
rect 292222 253058 292306 253294
rect 292542 253058 292574 253294
rect 291954 213614 292574 253058
rect 291954 213378 291986 213614
rect 292222 213378 292306 213614
rect 292542 213378 292574 213614
rect 291954 213294 292574 213378
rect 291954 213058 291986 213294
rect 292222 213058 292306 213294
rect 292542 213058 292574 213294
rect 291954 173614 292574 213058
rect 291954 173378 291986 173614
rect 292222 173378 292306 173614
rect 292542 173378 292574 173614
rect 291954 173294 292574 173378
rect 291954 173058 291986 173294
rect 292222 173058 292306 173294
rect 292542 173058 292574 173294
rect 291954 133614 292574 173058
rect 291954 133378 291986 133614
rect 292222 133378 292306 133614
rect 292542 133378 292574 133614
rect 291954 133294 292574 133378
rect 291954 133058 291986 133294
rect 292222 133058 292306 133294
rect 292542 133058 292574 133294
rect 291954 93614 292574 133058
rect 291954 93378 291986 93614
rect 292222 93378 292306 93614
rect 292542 93378 292574 93614
rect 291954 93294 292574 93378
rect 291954 93058 291986 93294
rect 292222 93058 292306 93294
rect 292542 93058 292574 93294
rect 291954 53614 292574 93058
rect 291954 53378 291986 53614
rect 292222 53378 292306 53614
rect 292542 53378 292574 53614
rect 291954 53294 292574 53378
rect 291954 53058 291986 53294
rect 292222 53058 292306 53294
rect 292542 53058 292574 53294
rect 291954 13614 292574 53058
rect 291954 13378 291986 13614
rect 292222 13378 292306 13614
rect 292542 13378 292574 13614
rect 291954 13294 292574 13378
rect 291954 13058 291986 13294
rect 292222 13058 292306 13294
rect 292542 13058 292574 13294
rect 271954 -7302 271986 -7066
rect 272222 -7302 272306 -7066
rect 272542 -7302 272574 -7066
rect 271954 -7386 272574 -7302
rect 271954 -7622 271986 -7386
rect 272222 -7622 272306 -7386
rect 272542 -7622 272574 -7386
rect 271954 -7654 272574 -7622
rect 291954 -6106 292574 13058
rect 293910 3365 293970 319363
rect 300794 302454 301414 341898
rect 304514 666174 305134 707162
rect 304514 665938 304546 666174
rect 304782 665938 304866 666174
rect 305102 665938 305134 666174
rect 304514 665854 305134 665938
rect 304514 665618 304546 665854
rect 304782 665618 304866 665854
rect 305102 665618 305134 665854
rect 304514 626174 305134 665618
rect 304514 625938 304546 626174
rect 304782 625938 304866 626174
rect 305102 625938 305134 626174
rect 304514 625854 305134 625938
rect 304514 625618 304546 625854
rect 304782 625618 304866 625854
rect 305102 625618 305134 625854
rect 304514 586174 305134 625618
rect 304514 585938 304546 586174
rect 304782 585938 304866 586174
rect 305102 585938 305134 586174
rect 304514 585854 305134 585938
rect 304514 585618 304546 585854
rect 304782 585618 304866 585854
rect 305102 585618 305134 585854
rect 304514 546174 305134 585618
rect 304514 545938 304546 546174
rect 304782 545938 304866 546174
rect 305102 545938 305134 546174
rect 304514 545854 305134 545938
rect 304514 545618 304546 545854
rect 304782 545618 304866 545854
rect 305102 545618 305134 545854
rect 304514 506174 305134 545618
rect 304514 505938 304546 506174
rect 304782 505938 304866 506174
rect 305102 505938 305134 506174
rect 304514 505854 305134 505938
rect 304514 505618 304546 505854
rect 304782 505618 304866 505854
rect 305102 505618 305134 505854
rect 304514 466174 305134 505618
rect 304514 465938 304546 466174
rect 304782 465938 304866 466174
rect 305102 465938 305134 466174
rect 304514 465854 305134 465938
rect 304514 465618 304546 465854
rect 304782 465618 304866 465854
rect 305102 465618 305134 465854
rect 304514 426174 305134 465618
rect 304514 425938 304546 426174
rect 304782 425938 304866 426174
rect 305102 425938 305134 426174
rect 304514 425854 305134 425938
rect 304514 425618 304546 425854
rect 304782 425618 304866 425854
rect 305102 425618 305134 425854
rect 304514 386174 305134 425618
rect 304514 385938 304546 386174
rect 304782 385938 304866 386174
rect 305102 385938 305134 386174
rect 304514 385854 305134 385938
rect 304514 385618 304546 385854
rect 304782 385618 304866 385854
rect 305102 385618 305134 385854
rect 304514 346174 305134 385618
rect 304514 345938 304546 346174
rect 304782 345938 304866 346174
rect 305102 345938 305134 346174
rect 304514 345854 305134 345938
rect 304514 345618 304546 345854
rect 304782 345618 304866 345854
rect 305102 345618 305134 345854
rect 303659 319428 303725 319429
rect 303659 319364 303660 319428
rect 303724 319364 303725 319428
rect 303659 319363 303725 319364
rect 300794 302218 300826 302454
rect 301382 302218 301414 302454
rect 300794 302134 301414 302218
rect 300794 301898 300826 302134
rect 301382 301898 301414 302134
rect 300794 262454 301414 301898
rect 300794 262218 300826 262454
rect 301382 262218 301414 262454
rect 300794 262134 301414 262218
rect 300794 261898 300826 262134
rect 301382 261898 301414 262134
rect 300794 222454 301414 261898
rect 300794 222218 300826 222454
rect 301382 222218 301414 222454
rect 300794 222134 301414 222218
rect 300794 221898 300826 222134
rect 301382 221898 301414 222134
rect 300794 182454 301414 221898
rect 300794 182218 300826 182454
rect 301382 182218 301414 182454
rect 300794 182134 301414 182218
rect 300794 181898 300826 182134
rect 301382 181898 301414 182134
rect 300794 142454 301414 181898
rect 300794 142218 300826 142454
rect 301382 142218 301414 142454
rect 300794 142134 301414 142218
rect 300794 141898 300826 142134
rect 301382 141898 301414 142134
rect 300794 102454 301414 141898
rect 300794 102218 300826 102454
rect 301062 102218 301146 102454
rect 301382 102218 301414 102454
rect 300794 102134 301414 102218
rect 300794 101898 300826 102134
rect 301062 101898 301146 102134
rect 301382 101898 301414 102134
rect 300794 62454 301414 101898
rect 300794 62218 300826 62454
rect 301062 62218 301146 62454
rect 301382 62218 301414 62454
rect 300794 62134 301414 62218
rect 300794 61898 300826 62134
rect 301062 61898 301146 62134
rect 301382 61898 301414 62134
rect 300794 22454 301414 61898
rect 300794 22218 300826 22454
rect 301062 22218 301146 22454
rect 301382 22218 301414 22454
rect 300794 22134 301414 22218
rect 300794 21898 300826 22134
rect 301062 21898 301146 22134
rect 301382 21898 301414 22134
rect 293907 3364 293973 3365
rect 293907 3300 293908 3364
rect 293972 3300 293973 3364
rect 293907 3299 293973 3300
rect 300794 -1306 301414 21898
rect 303662 3909 303722 319363
rect 304514 306174 305134 345618
rect 304514 305938 304546 306174
rect 304782 305938 304866 306174
rect 305102 305938 305134 306174
rect 304514 305854 305134 305938
rect 304514 305618 304546 305854
rect 304782 305618 304866 305854
rect 305102 305618 305134 305854
rect 304514 266174 305134 305618
rect 304514 265938 304546 266174
rect 304782 265938 304866 266174
rect 305102 265938 305134 266174
rect 304514 265854 305134 265938
rect 304514 265618 304546 265854
rect 304782 265618 304866 265854
rect 305102 265618 305134 265854
rect 304514 226174 305134 265618
rect 304514 225938 304546 226174
rect 304782 225938 304866 226174
rect 305102 225938 305134 226174
rect 304514 225854 305134 225938
rect 304514 225618 304546 225854
rect 304782 225618 304866 225854
rect 305102 225618 305134 225854
rect 304514 186174 305134 225618
rect 304514 185938 304546 186174
rect 304782 185938 304866 186174
rect 305102 185938 305134 186174
rect 304514 185854 305134 185938
rect 304514 185618 304546 185854
rect 304782 185618 304866 185854
rect 305102 185618 305134 185854
rect 304514 146174 305134 185618
rect 304514 145938 304546 146174
rect 304782 145938 304866 146174
rect 305102 145938 305134 146174
rect 304514 145854 305134 145938
rect 304514 145618 304546 145854
rect 304782 145618 304866 145854
rect 305102 145618 305134 145854
rect 304514 106174 305134 145618
rect 304514 105938 304546 106174
rect 304782 105938 304866 106174
rect 305102 105938 305134 106174
rect 304514 105854 305134 105938
rect 304514 105618 304546 105854
rect 304782 105618 304866 105854
rect 305102 105618 305134 105854
rect 304514 66174 305134 105618
rect 304514 65938 304546 66174
rect 304782 65938 304866 66174
rect 305102 65938 305134 66174
rect 304514 65854 305134 65938
rect 304514 65618 304546 65854
rect 304782 65618 304866 65854
rect 305102 65618 305134 65854
rect 304514 26174 305134 65618
rect 304514 25938 304546 26174
rect 304782 25938 304866 26174
rect 305102 25938 305134 26174
rect 304514 25854 305134 25938
rect 304514 25618 304546 25854
rect 304782 25618 304866 25854
rect 305102 25618 305134 25854
rect 303659 3908 303725 3909
rect 303659 3844 303660 3908
rect 303724 3844 303725 3908
rect 303659 3843 303725 3844
rect 300794 -1542 300826 -1306
rect 301062 -1542 301146 -1306
rect 301382 -1542 301414 -1306
rect 300794 -1626 301414 -1542
rect 300794 -1862 300826 -1626
rect 301062 -1862 301146 -1626
rect 301382 -1862 301414 -1626
rect 300794 -1894 301414 -1862
rect 304514 -3226 305134 25618
rect 304514 -3462 304546 -3226
rect 304782 -3462 304866 -3226
rect 305102 -3462 305134 -3226
rect 304514 -3546 305134 -3462
rect 304514 -3782 304546 -3546
rect 304782 -3782 304866 -3546
rect 305102 -3782 305134 -3546
rect 304514 -3814 305134 -3782
rect 308234 669894 308854 709082
rect 308234 669658 308266 669894
rect 308502 669658 308586 669894
rect 308822 669658 308854 669894
rect 308234 669574 308854 669658
rect 308234 669338 308266 669574
rect 308502 669338 308586 669574
rect 308822 669338 308854 669574
rect 308234 629894 308854 669338
rect 308234 629658 308266 629894
rect 308502 629658 308586 629894
rect 308822 629658 308854 629894
rect 308234 629574 308854 629658
rect 308234 629338 308266 629574
rect 308502 629338 308586 629574
rect 308822 629338 308854 629574
rect 308234 589894 308854 629338
rect 308234 589658 308266 589894
rect 308502 589658 308586 589894
rect 308822 589658 308854 589894
rect 308234 589574 308854 589658
rect 308234 589338 308266 589574
rect 308502 589338 308586 589574
rect 308822 589338 308854 589574
rect 308234 549894 308854 589338
rect 308234 549658 308266 549894
rect 308502 549658 308586 549894
rect 308822 549658 308854 549894
rect 308234 549574 308854 549658
rect 308234 549338 308266 549574
rect 308502 549338 308586 549574
rect 308822 549338 308854 549574
rect 308234 509894 308854 549338
rect 308234 509658 308266 509894
rect 308502 509658 308586 509894
rect 308822 509658 308854 509894
rect 308234 509574 308854 509658
rect 308234 509338 308266 509574
rect 308502 509338 308586 509574
rect 308822 509338 308854 509574
rect 308234 469894 308854 509338
rect 308234 469658 308266 469894
rect 308502 469658 308586 469894
rect 308822 469658 308854 469894
rect 308234 469574 308854 469658
rect 308234 469338 308266 469574
rect 308502 469338 308586 469574
rect 308822 469338 308854 469574
rect 308234 429894 308854 469338
rect 308234 429658 308266 429894
rect 308502 429658 308586 429894
rect 308822 429658 308854 429894
rect 308234 429574 308854 429658
rect 308234 429338 308266 429574
rect 308502 429338 308586 429574
rect 308822 429338 308854 429574
rect 308234 389894 308854 429338
rect 308234 389658 308266 389894
rect 308502 389658 308586 389894
rect 308822 389658 308854 389894
rect 308234 389574 308854 389658
rect 308234 389338 308266 389574
rect 308502 389338 308586 389574
rect 308822 389338 308854 389574
rect 308234 349894 308854 389338
rect 308234 349658 308266 349894
rect 308502 349658 308586 349894
rect 308822 349658 308854 349894
rect 308234 349574 308854 349658
rect 308234 349338 308266 349574
rect 308502 349338 308586 349574
rect 308822 349338 308854 349574
rect 308234 309894 308854 349338
rect 308234 309658 308266 309894
rect 308502 309658 308586 309894
rect 308822 309658 308854 309894
rect 308234 309574 308854 309658
rect 308234 309338 308266 309574
rect 308502 309338 308586 309574
rect 308822 309338 308854 309574
rect 308234 269894 308854 309338
rect 308234 269658 308266 269894
rect 308502 269658 308586 269894
rect 308822 269658 308854 269894
rect 308234 269574 308854 269658
rect 308234 269338 308266 269574
rect 308502 269338 308586 269574
rect 308822 269338 308854 269574
rect 308234 229894 308854 269338
rect 308234 229658 308266 229894
rect 308502 229658 308586 229894
rect 308822 229658 308854 229894
rect 308234 229574 308854 229658
rect 308234 229338 308266 229574
rect 308502 229338 308586 229574
rect 308822 229338 308854 229574
rect 308234 189894 308854 229338
rect 308234 189658 308266 189894
rect 308502 189658 308586 189894
rect 308822 189658 308854 189894
rect 308234 189574 308854 189658
rect 308234 189338 308266 189574
rect 308502 189338 308586 189574
rect 308822 189338 308854 189574
rect 308234 149894 308854 189338
rect 308234 149658 308266 149894
rect 308502 149658 308586 149894
rect 308822 149658 308854 149894
rect 308234 149574 308854 149658
rect 308234 149338 308266 149574
rect 308502 149338 308586 149574
rect 308822 149338 308854 149574
rect 308234 109894 308854 149338
rect 308234 109658 308266 109894
rect 308502 109658 308586 109894
rect 308822 109658 308854 109894
rect 308234 109574 308854 109658
rect 308234 109338 308266 109574
rect 308502 109338 308586 109574
rect 308822 109338 308854 109574
rect 308234 69894 308854 109338
rect 308234 69658 308266 69894
rect 308502 69658 308586 69894
rect 308822 69658 308854 69894
rect 308234 69574 308854 69658
rect 308234 69338 308266 69574
rect 308502 69338 308586 69574
rect 308822 69338 308854 69574
rect 308234 29894 308854 69338
rect 308234 29658 308266 29894
rect 308502 29658 308586 29894
rect 308822 29658 308854 29894
rect 308234 29574 308854 29658
rect 308234 29338 308266 29574
rect 308502 29338 308586 29574
rect 308822 29338 308854 29574
rect 308234 -5146 308854 29338
rect 308234 -5382 308266 -5146
rect 308502 -5382 308586 -5146
rect 308822 -5382 308854 -5146
rect 308234 -5466 308854 -5382
rect 308234 -5702 308266 -5466
rect 308502 -5702 308586 -5466
rect 308822 -5702 308854 -5466
rect 308234 -5734 308854 -5702
rect 311954 673614 312574 711002
rect 331954 710598 332574 711590
rect 331954 710362 331986 710598
rect 332222 710362 332306 710598
rect 332542 710362 332574 710598
rect 331954 710278 332574 710362
rect 331954 710042 331986 710278
rect 332222 710042 332306 710278
rect 332542 710042 332574 710278
rect 328234 708678 328854 709670
rect 328234 708442 328266 708678
rect 328502 708442 328586 708678
rect 328822 708442 328854 708678
rect 328234 708358 328854 708442
rect 328234 708122 328266 708358
rect 328502 708122 328586 708358
rect 328822 708122 328854 708358
rect 324514 706758 325134 707750
rect 324514 706522 324546 706758
rect 324782 706522 324866 706758
rect 325102 706522 325134 706758
rect 324514 706438 325134 706522
rect 324514 706202 324546 706438
rect 324782 706202 324866 706438
rect 325102 706202 325134 706438
rect 311954 673378 311986 673614
rect 312222 673378 312306 673614
rect 312542 673378 312574 673614
rect 311954 673294 312574 673378
rect 311954 673058 311986 673294
rect 312222 673058 312306 673294
rect 312542 673058 312574 673294
rect 311954 633614 312574 673058
rect 311954 633378 311986 633614
rect 312222 633378 312306 633614
rect 312542 633378 312574 633614
rect 311954 633294 312574 633378
rect 311954 633058 311986 633294
rect 312222 633058 312306 633294
rect 312542 633058 312574 633294
rect 311954 593614 312574 633058
rect 311954 593378 311986 593614
rect 312222 593378 312306 593614
rect 312542 593378 312574 593614
rect 311954 593294 312574 593378
rect 311954 593058 311986 593294
rect 312222 593058 312306 593294
rect 312542 593058 312574 593294
rect 311954 553614 312574 593058
rect 311954 553378 311986 553614
rect 312222 553378 312306 553614
rect 312542 553378 312574 553614
rect 311954 553294 312574 553378
rect 311954 553058 311986 553294
rect 312222 553058 312306 553294
rect 312542 553058 312574 553294
rect 311954 513614 312574 553058
rect 311954 513378 311986 513614
rect 312222 513378 312306 513614
rect 312542 513378 312574 513614
rect 311954 513294 312574 513378
rect 311954 513058 311986 513294
rect 312222 513058 312306 513294
rect 312542 513058 312574 513294
rect 311954 473614 312574 513058
rect 311954 473378 311986 473614
rect 312222 473378 312306 473614
rect 312542 473378 312574 473614
rect 311954 473294 312574 473378
rect 311954 473058 311986 473294
rect 312222 473058 312306 473294
rect 312542 473058 312574 473294
rect 311954 433614 312574 473058
rect 311954 433378 311986 433614
rect 312222 433378 312306 433614
rect 312542 433378 312574 433614
rect 311954 433294 312574 433378
rect 311954 433058 311986 433294
rect 312222 433058 312306 433294
rect 312542 433058 312574 433294
rect 311954 393614 312574 433058
rect 311954 393378 311986 393614
rect 312222 393378 312306 393614
rect 312542 393378 312574 393614
rect 311954 393294 312574 393378
rect 311954 393058 311986 393294
rect 312222 393058 312306 393294
rect 312542 393058 312574 393294
rect 311954 353614 312574 393058
rect 311954 353378 311986 353614
rect 312222 353378 312306 353614
rect 312542 353378 312574 353614
rect 311954 353294 312574 353378
rect 311954 353058 311986 353294
rect 312222 353058 312306 353294
rect 312542 353058 312574 353294
rect 311954 313614 312574 353058
rect 320794 704838 321414 705830
rect 320794 704602 320826 704838
rect 321062 704602 321146 704838
rect 321382 704602 321414 704838
rect 320794 704518 321414 704602
rect 320794 704282 320826 704518
rect 321062 704282 321146 704518
rect 321382 704282 321414 704518
rect 320794 682454 321414 704282
rect 320794 682218 320826 682454
rect 321062 682218 321146 682454
rect 321382 682218 321414 682454
rect 320794 682134 321414 682218
rect 320794 681898 320826 682134
rect 321062 681898 321146 682134
rect 321382 681898 321414 682134
rect 320794 642454 321414 681898
rect 320794 642218 320826 642454
rect 321062 642218 321146 642454
rect 321382 642218 321414 642454
rect 320794 642134 321414 642218
rect 320794 641898 320826 642134
rect 321062 641898 321146 642134
rect 321382 641898 321414 642134
rect 320794 602454 321414 641898
rect 320794 602218 320826 602454
rect 321062 602218 321146 602454
rect 321382 602218 321414 602454
rect 320794 602134 321414 602218
rect 320794 601898 320826 602134
rect 321062 601898 321146 602134
rect 321382 601898 321414 602134
rect 320794 562454 321414 601898
rect 320794 562218 320826 562454
rect 321062 562218 321146 562454
rect 321382 562218 321414 562454
rect 320794 562134 321414 562218
rect 320794 561898 320826 562134
rect 321062 561898 321146 562134
rect 321382 561898 321414 562134
rect 320794 522454 321414 561898
rect 320794 522218 320826 522454
rect 321062 522218 321146 522454
rect 321382 522218 321414 522454
rect 320794 522134 321414 522218
rect 320794 521898 320826 522134
rect 321062 521898 321146 522134
rect 321382 521898 321414 522134
rect 320794 482454 321414 521898
rect 320794 482218 320826 482454
rect 321062 482218 321146 482454
rect 321382 482218 321414 482454
rect 320794 482134 321414 482218
rect 320794 481898 320826 482134
rect 321062 481898 321146 482134
rect 321382 481898 321414 482134
rect 320794 442454 321414 481898
rect 320794 442218 320826 442454
rect 321062 442218 321146 442454
rect 321382 442218 321414 442454
rect 320794 442134 321414 442218
rect 320794 441898 320826 442134
rect 321062 441898 321146 442134
rect 321382 441898 321414 442134
rect 320794 402454 321414 441898
rect 320794 402218 320826 402454
rect 321062 402218 321146 402454
rect 321382 402218 321414 402454
rect 320794 402134 321414 402218
rect 320794 401898 320826 402134
rect 321062 401898 321146 402134
rect 321382 401898 321414 402134
rect 320794 362454 321414 401898
rect 320794 362218 320826 362454
rect 321062 362218 321146 362454
rect 321382 362218 321414 362454
rect 320794 362134 321414 362218
rect 320794 361898 320826 362134
rect 321062 361898 321146 362134
rect 321382 361898 321414 362134
rect 320794 322454 321414 361898
rect 320794 322218 320826 322454
rect 321062 322218 321146 322454
rect 321382 322218 321414 322454
rect 320794 322134 321414 322218
rect 320794 321898 320826 322134
rect 321062 321898 321146 322134
rect 321382 321898 321414 322134
rect 314699 319428 314765 319429
rect 314699 319364 314700 319428
rect 314764 319364 314765 319428
rect 314699 319363 314765 319364
rect 311954 313378 311986 313614
rect 312222 313378 312306 313614
rect 312542 313378 312574 313614
rect 311954 313294 312574 313378
rect 311954 313058 311986 313294
rect 312222 313058 312306 313294
rect 312542 313058 312574 313294
rect 311954 273614 312574 313058
rect 311954 273378 311986 273614
rect 312222 273378 312306 273614
rect 312542 273378 312574 273614
rect 311954 273294 312574 273378
rect 311954 273058 311986 273294
rect 312222 273058 312306 273294
rect 312542 273058 312574 273294
rect 311954 233614 312574 273058
rect 311954 233378 311986 233614
rect 312222 233378 312306 233614
rect 312542 233378 312574 233614
rect 311954 233294 312574 233378
rect 311954 233058 311986 233294
rect 312222 233058 312306 233294
rect 312542 233058 312574 233294
rect 311954 193614 312574 233058
rect 311954 193378 311986 193614
rect 312222 193378 312306 193614
rect 312542 193378 312574 193614
rect 311954 193294 312574 193378
rect 311954 193058 311986 193294
rect 312222 193058 312306 193294
rect 312542 193058 312574 193294
rect 311954 153614 312574 193058
rect 311954 153378 311986 153614
rect 312222 153378 312306 153614
rect 312542 153378 312574 153614
rect 311954 153294 312574 153378
rect 311954 153058 311986 153294
rect 312222 153058 312306 153294
rect 312542 153058 312574 153294
rect 311954 113614 312574 153058
rect 311954 113378 311986 113614
rect 312222 113378 312306 113614
rect 312542 113378 312574 113614
rect 311954 113294 312574 113378
rect 311954 113058 311986 113294
rect 312222 113058 312306 113294
rect 312542 113058 312574 113294
rect 311954 73614 312574 113058
rect 311954 73378 311986 73614
rect 312222 73378 312306 73614
rect 312542 73378 312574 73614
rect 311954 73294 312574 73378
rect 311954 73058 311986 73294
rect 312222 73058 312306 73294
rect 312542 73058 312574 73294
rect 311954 33614 312574 73058
rect 311954 33378 311986 33614
rect 312222 33378 312306 33614
rect 312542 33378 312574 33614
rect 311954 33294 312574 33378
rect 311954 33058 311986 33294
rect 312222 33058 312306 33294
rect 312542 33058 312574 33294
rect 291954 -6342 291986 -6106
rect 292222 -6342 292306 -6106
rect 292542 -6342 292574 -6106
rect 291954 -6426 292574 -6342
rect 291954 -6662 291986 -6426
rect 292222 -6662 292306 -6426
rect 292542 -6662 292574 -6426
rect 291954 -7654 292574 -6662
rect 311954 -7066 312574 33058
rect 314702 3637 314762 319363
rect 320794 282454 321414 321898
rect 320794 282218 320826 282454
rect 321062 282218 321146 282454
rect 321382 282218 321414 282454
rect 320794 282134 321414 282218
rect 320794 281898 320826 282134
rect 321062 281898 321146 282134
rect 321382 281898 321414 282134
rect 320794 242454 321414 281898
rect 320794 242218 320826 242454
rect 321062 242218 321146 242454
rect 321382 242218 321414 242454
rect 320794 242134 321414 242218
rect 320794 241898 320826 242134
rect 321062 241898 321146 242134
rect 321382 241898 321414 242134
rect 320794 202454 321414 241898
rect 320794 202218 320826 202454
rect 321062 202218 321146 202454
rect 321382 202218 321414 202454
rect 320794 202134 321414 202218
rect 320794 201898 320826 202134
rect 321062 201898 321146 202134
rect 321382 201898 321414 202134
rect 320794 162454 321414 201898
rect 320794 162218 320826 162454
rect 321062 162218 321146 162454
rect 321382 162218 321414 162454
rect 320794 162134 321414 162218
rect 320794 161898 320826 162134
rect 321062 161898 321146 162134
rect 321382 161898 321414 162134
rect 320794 122454 321414 161898
rect 320794 122218 320826 122454
rect 321062 122218 321146 122454
rect 321382 122218 321414 122454
rect 320794 122134 321414 122218
rect 320794 121898 320826 122134
rect 321062 121898 321146 122134
rect 321382 121898 321414 122134
rect 320794 82454 321414 121898
rect 320794 82218 320826 82454
rect 321062 82218 321146 82454
rect 321382 82218 321414 82454
rect 320794 82134 321414 82218
rect 320794 81898 320826 82134
rect 321062 81898 321146 82134
rect 321382 81898 321414 82134
rect 320794 42454 321414 81898
rect 320794 42218 320826 42454
rect 321062 42218 321146 42454
rect 321382 42218 321414 42454
rect 320794 42134 321414 42218
rect 320794 41898 320826 42134
rect 321062 41898 321146 42134
rect 321382 41898 321414 42134
rect 314699 3636 314765 3637
rect 314699 3572 314700 3636
rect 314764 3572 314765 3636
rect 314699 3571 314765 3572
rect 320794 2454 321414 41898
rect 320794 2218 320826 2454
rect 321062 2218 321146 2454
rect 321382 2218 321414 2454
rect 320794 2134 321414 2218
rect 320794 1898 320826 2134
rect 321062 1898 321146 2134
rect 321382 1898 321414 2134
rect 320794 -346 321414 1898
rect 320794 -582 320826 -346
rect 321062 -582 321146 -346
rect 321382 -582 321414 -346
rect 320794 -666 321414 -582
rect 320794 -902 320826 -666
rect 321062 -902 321146 -666
rect 321382 -902 321414 -666
rect 320794 -1894 321414 -902
rect 324514 686174 325134 706202
rect 324514 685938 324546 686174
rect 324782 685938 324866 686174
rect 325102 685938 325134 686174
rect 324514 685854 325134 685938
rect 324514 685618 324546 685854
rect 324782 685618 324866 685854
rect 325102 685618 325134 685854
rect 324514 646174 325134 685618
rect 324514 645938 324546 646174
rect 324782 645938 324866 646174
rect 325102 645938 325134 646174
rect 324514 645854 325134 645938
rect 324514 645618 324546 645854
rect 324782 645618 324866 645854
rect 325102 645618 325134 645854
rect 324514 606174 325134 645618
rect 324514 605938 324546 606174
rect 324782 605938 324866 606174
rect 325102 605938 325134 606174
rect 324514 605854 325134 605938
rect 324514 605618 324546 605854
rect 324782 605618 324866 605854
rect 325102 605618 325134 605854
rect 324514 566174 325134 605618
rect 324514 565938 324546 566174
rect 324782 565938 324866 566174
rect 325102 565938 325134 566174
rect 324514 565854 325134 565938
rect 324514 565618 324546 565854
rect 324782 565618 324866 565854
rect 325102 565618 325134 565854
rect 324514 526174 325134 565618
rect 324514 525938 324546 526174
rect 324782 525938 324866 526174
rect 325102 525938 325134 526174
rect 324514 525854 325134 525938
rect 324514 525618 324546 525854
rect 324782 525618 324866 525854
rect 325102 525618 325134 525854
rect 324514 486174 325134 525618
rect 324514 485938 324546 486174
rect 324782 485938 324866 486174
rect 325102 485938 325134 486174
rect 324514 485854 325134 485938
rect 324514 485618 324546 485854
rect 324782 485618 324866 485854
rect 325102 485618 325134 485854
rect 324514 446174 325134 485618
rect 324514 445938 324546 446174
rect 324782 445938 324866 446174
rect 325102 445938 325134 446174
rect 324514 445854 325134 445938
rect 324514 445618 324546 445854
rect 324782 445618 324866 445854
rect 325102 445618 325134 445854
rect 324514 406174 325134 445618
rect 324514 405938 324546 406174
rect 324782 405938 324866 406174
rect 325102 405938 325134 406174
rect 324514 405854 325134 405938
rect 324514 405618 324546 405854
rect 324782 405618 324866 405854
rect 325102 405618 325134 405854
rect 324514 366174 325134 405618
rect 324514 365938 324546 366174
rect 324782 365938 324866 366174
rect 325102 365938 325134 366174
rect 324514 365854 325134 365938
rect 324514 365618 324546 365854
rect 324782 365618 324866 365854
rect 325102 365618 325134 365854
rect 324514 326174 325134 365618
rect 324514 325938 324546 326174
rect 324782 325938 324866 326174
rect 325102 325938 325134 326174
rect 324514 325854 325134 325938
rect 324514 325618 324546 325854
rect 324782 325618 324866 325854
rect 325102 325618 325134 325854
rect 324514 286174 325134 325618
rect 324514 285938 324546 286174
rect 324782 285938 324866 286174
rect 325102 285938 325134 286174
rect 324514 285854 325134 285938
rect 324514 285618 324546 285854
rect 324782 285618 324866 285854
rect 325102 285618 325134 285854
rect 324514 246174 325134 285618
rect 324514 245938 324546 246174
rect 324782 245938 324866 246174
rect 325102 245938 325134 246174
rect 324514 245854 325134 245938
rect 324514 245618 324546 245854
rect 324782 245618 324866 245854
rect 325102 245618 325134 245854
rect 324514 206174 325134 245618
rect 324514 205938 324546 206174
rect 324782 205938 324866 206174
rect 325102 205938 325134 206174
rect 324514 205854 325134 205938
rect 324514 205618 324546 205854
rect 324782 205618 324866 205854
rect 325102 205618 325134 205854
rect 324514 166174 325134 205618
rect 324514 165938 324546 166174
rect 324782 165938 324866 166174
rect 325102 165938 325134 166174
rect 324514 165854 325134 165938
rect 324514 165618 324546 165854
rect 324782 165618 324866 165854
rect 325102 165618 325134 165854
rect 324514 126174 325134 165618
rect 324514 125938 324546 126174
rect 324782 125938 324866 126174
rect 325102 125938 325134 126174
rect 324514 125854 325134 125938
rect 324514 125618 324546 125854
rect 324782 125618 324866 125854
rect 325102 125618 325134 125854
rect 324514 86174 325134 125618
rect 324514 85938 324546 86174
rect 324782 85938 324866 86174
rect 325102 85938 325134 86174
rect 324514 85854 325134 85938
rect 324514 85618 324546 85854
rect 324782 85618 324866 85854
rect 325102 85618 325134 85854
rect 324514 46174 325134 85618
rect 324514 45938 324546 46174
rect 324782 45938 324866 46174
rect 325102 45938 325134 46174
rect 324514 45854 325134 45938
rect 324514 45618 324546 45854
rect 324782 45618 324866 45854
rect 325102 45618 325134 45854
rect 324514 6174 325134 45618
rect 324514 5938 324546 6174
rect 324782 5938 324866 6174
rect 325102 5938 325134 6174
rect 324514 5854 325134 5938
rect 324514 5618 324546 5854
rect 324782 5618 324866 5854
rect 325102 5618 325134 5854
rect 324514 -2266 325134 5618
rect 324514 -2502 324546 -2266
rect 324782 -2502 324866 -2266
rect 325102 -2502 325134 -2266
rect 324514 -2586 325134 -2502
rect 324514 -2822 324546 -2586
rect 324782 -2822 324866 -2586
rect 325102 -2822 325134 -2586
rect 324514 -3814 325134 -2822
rect 328234 689894 328854 708122
rect 328234 689658 328266 689894
rect 328502 689658 328586 689894
rect 328822 689658 328854 689894
rect 328234 689574 328854 689658
rect 328234 689338 328266 689574
rect 328502 689338 328586 689574
rect 328822 689338 328854 689574
rect 328234 649894 328854 689338
rect 328234 649658 328266 649894
rect 328502 649658 328586 649894
rect 328822 649658 328854 649894
rect 328234 649574 328854 649658
rect 328234 649338 328266 649574
rect 328502 649338 328586 649574
rect 328822 649338 328854 649574
rect 328234 609894 328854 649338
rect 328234 609658 328266 609894
rect 328502 609658 328586 609894
rect 328822 609658 328854 609894
rect 328234 609574 328854 609658
rect 328234 609338 328266 609574
rect 328502 609338 328586 609574
rect 328822 609338 328854 609574
rect 328234 569894 328854 609338
rect 328234 569658 328266 569894
rect 328502 569658 328586 569894
rect 328822 569658 328854 569894
rect 328234 569574 328854 569658
rect 328234 569338 328266 569574
rect 328502 569338 328586 569574
rect 328822 569338 328854 569574
rect 328234 529894 328854 569338
rect 328234 529658 328266 529894
rect 328502 529658 328586 529894
rect 328822 529658 328854 529894
rect 328234 529574 328854 529658
rect 328234 529338 328266 529574
rect 328502 529338 328586 529574
rect 328822 529338 328854 529574
rect 328234 489894 328854 529338
rect 328234 489658 328266 489894
rect 328502 489658 328586 489894
rect 328822 489658 328854 489894
rect 328234 489574 328854 489658
rect 328234 489338 328266 489574
rect 328502 489338 328586 489574
rect 328822 489338 328854 489574
rect 328234 449894 328854 489338
rect 328234 449658 328266 449894
rect 328502 449658 328586 449894
rect 328822 449658 328854 449894
rect 328234 449574 328854 449658
rect 328234 449338 328266 449574
rect 328502 449338 328586 449574
rect 328822 449338 328854 449574
rect 328234 409894 328854 449338
rect 328234 409658 328266 409894
rect 328502 409658 328586 409894
rect 328822 409658 328854 409894
rect 328234 409574 328854 409658
rect 328234 409338 328266 409574
rect 328502 409338 328586 409574
rect 328822 409338 328854 409574
rect 328234 369894 328854 409338
rect 328234 369658 328266 369894
rect 328502 369658 328586 369894
rect 328822 369658 328854 369894
rect 328234 369574 328854 369658
rect 328234 369338 328266 369574
rect 328502 369338 328586 369574
rect 328822 369338 328854 369574
rect 328234 329894 328854 369338
rect 328234 329658 328266 329894
rect 328502 329658 328586 329894
rect 328822 329658 328854 329894
rect 328234 329574 328854 329658
rect 328234 329338 328266 329574
rect 328502 329338 328586 329574
rect 328822 329338 328854 329574
rect 328234 289894 328854 329338
rect 328234 289658 328266 289894
rect 328502 289658 328586 289894
rect 328822 289658 328854 289894
rect 328234 289574 328854 289658
rect 328234 289338 328266 289574
rect 328502 289338 328586 289574
rect 328822 289338 328854 289574
rect 328234 249894 328854 289338
rect 328234 249658 328266 249894
rect 328502 249658 328586 249894
rect 328822 249658 328854 249894
rect 328234 249574 328854 249658
rect 328234 249338 328266 249574
rect 328502 249338 328586 249574
rect 328822 249338 328854 249574
rect 328234 209894 328854 249338
rect 328234 209658 328266 209894
rect 328502 209658 328586 209894
rect 328822 209658 328854 209894
rect 328234 209574 328854 209658
rect 328234 209338 328266 209574
rect 328502 209338 328586 209574
rect 328822 209338 328854 209574
rect 328234 169894 328854 209338
rect 328234 169658 328266 169894
rect 328502 169658 328586 169894
rect 328822 169658 328854 169894
rect 328234 169574 328854 169658
rect 328234 169338 328266 169574
rect 328502 169338 328586 169574
rect 328822 169338 328854 169574
rect 328234 129894 328854 169338
rect 328234 129658 328266 129894
rect 328502 129658 328586 129894
rect 328822 129658 328854 129894
rect 328234 129574 328854 129658
rect 328234 129338 328266 129574
rect 328502 129338 328586 129574
rect 328822 129338 328854 129574
rect 328234 89894 328854 129338
rect 328234 89658 328266 89894
rect 328502 89658 328586 89894
rect 328822 89658 328854 89894
rect 328234 89574 328854 89658
rect 328234 89338 328266 89574
rect 328502 89338 328586 89574
rect 328822 89338 328854 89574
rect 328234 49894 328854 89338
rect 328234 49658 328266 49894
rect 328502 49658 328586 49894
rect 328822 49658 328854 49894
rect 328234 49574 328854 49658
rect 328234 49338 328266 49574
rect 328502 49338 328586 49574
rect 328822 49338 328854 49574
rect 328234 9894 328854 49338
rect 328234 9658 328266 9894
rect 328502 9658 328586 9894
rect 328822 9658 328854 9894
rect 328234 9574 328854 9658
rect 328234 9338 328266 9574
rect 328502 9338 328586 9574
rect 328822 9338 328854 9574
rect 328234 -4186 328854 9338
rect 328234 -4422 328266 -4186
rect 328502 -4422 328586 -4186
rect 328822 -4422 328854 -4186
rect 328234 -4506 328854 -4422
rect 328234 -4742 328266 -4506
rect 328502 -4742 328586 -4506
rect 328822 -4742 328854 -4506
rect 328234 -5734 328854 -4742
rect 331954 693614 332574 710042
rect 351954 711558 352574 711590
rect 351954 711322 351986 711558
rect 352222 711322 352306 711558
rect 352542 711322 352574 711558
rect 351954 711238 352574 711322
rect 351954 711002 351986 711238
rect 352222 711002 352306 711238
rect 352542 711002 352574 711238
rect 348234 709638 348854 709670
rect 348234 709402 348266 709638
rect 348502 709402 348586 709638
rect 348822 709402 348854 709638
rect 348234 709318 348854 709402
rect 348234 709082 348266 709318
rect 348502 709082 348586 709318
rect 348822 709082 348854 709318
rect 344514 707718 345134 707750
rect 344514 707482 344546 707718
rect 344782 707482 344866 707718
rect 345102 707482 345134 707718
rect 344514 707398 345134 707482
rect 344514 707162 344546 707398
rect 344782 707162 344866 707398
rect 345102 707162 345134 707398
rect 331954 693378 331986 693614
rect 332222 693378 332306 693614
rect 332542 693378 332574 693614
rect 331954 693294 332574 693378
rect 331954 693058 331986 693294
rect 332222 693058 332306 693294
rect 332542 693058 332574 693294
rect 331954 653614 332574 693058
rect 331954 653378 331986 653614
rect 332222 653378 332306 653614
rect 332542 653378 332574 653614
rect 331954 653294 332574 653378
rect 331954 653058 331986 653294
rect 332222 653058 332306 653294
rect 332542 653058 332574 653294
rect 331954 613614 332574 653058
rect 331954 613378 331986 613614
rect 332222 613378 332306 613614
rect 332542 613378 332574 613614
rect 331954 613294 332574 613378
rect 331954 613058 331986 613294
rect 332222 613058 332306 613294
rect 332542 613058 332574 613294
rect 331954 573614 332574 613058
rect 331954 573378 331986 573614
rect 332222 573378 332306 573614
rect 332542 573378 332574 573614
rect 331954 573294 332574 573378
rect 331954 573058 331986 573294
rect 332222 573058 332306 573294
rect 332542 573058 332574 573294
rect 331954 533614 332574 573058
rect 331954 533378 331986 533614
rect 332222 533378 332306 533614
rect 332542 533378 332574 533614
rect 331954 533294 332574 533378
rect 331954 533058 331986 533294
rect 332222 533058 332306 533294
rect 332542 533058 332574 533294
rect 331954 493614 332574 533058
rect 331954 493378 331986 493614
rect 332222 493378 332306 493614
rect 332542 493378 332574 493614
rect 331954 493294 332574 493378
rect 331954 493058 331986 493294
rect 332222 493058 332306 493294
rect 332542 493058 332574 493294
rect 331954 453614 332574 493058
rect 331954 453378 331986 453614
rect 332222 453378 332306 453614
rect 332542 453378 332574 453614
rect 331954 453294 332574 453378
rect 331954 453058 331986 453294
rect 332222 453058 332306 453294
rect 332542 453058 332574 453294
rect 331954 413614 332574 453058
rect 331954 413378 331986 413614
rect 332222 413378 332306 413614
rect 332542 413378 332574 413614
rect 331954 413294 332574 413378
rect 331954 413058 331986 413294
rect 332222 413058 332306 413294
rect 332542 413058 332574 413294
rect 331954 373614 332574 413058
rect 331954 373378 331986 373614
rect 332222 373378 332306 373614
rect 332542 373378 332574 373614
rect 331954 373294 332574 373378
rect 331954 373058 331986 373294
rect 332222 373058 332306 373294
rect 332542 373058 332574 373294
rect 331954 333614 332574 373058
rect 331954 333378 331986 333614
rect 332222 333378 332306 333614
rect 332542 333378 332574 333614
rect 331954 333294 332574 333378
rect 331954 333058 331986 333294
rect 332222 333058 332306 333294
rect 332542 333058 332574 333294
rect 331954 293614 332574 333058
rect 331954 293378 331986 293614
rect 332222 293378 332306 293614
rect 332542 293378 332574 293614
rect 331954 293294 332574 293378
rect 331954 293058 331986 293294
rect 332222 293058 332306 293294
rect 332542 293058 332574 293294
rect 331954 253614 332574 293058
rect 331954 253378 331986 253614
rect 332222 253378 332306 253614
rect 332542 253378 332574 253614
rect 331954 253294 332574 253378
rect 331954 253058 331986 253294
rect 332222 253058 332306 253294
rect 332542 253058 332574 253294
rect 331954 213614 332574 253058
rect 331954 213378 331986 213614
rect 332222 213378 332306 213614
rect 332542 213378 332574 213614
rect 331954 213294 332574 213378
rect 331954 213058 331986 213294
rect 332222 213058 332306 213294
rect 332542 213058 332574 213294
rect 331954 173614 332574 213058
rect 331954 173378 331986 173614
rect 332222 173378 332306 173614
rect 332542 173378 332574 173614
rect 331954 173294 332574 173378
rect 331954 173058 331986 173294
rect 332222 173058 332306 173294
rect 332542 173058 332574 173294
rect 331954 133614 332574 173058
rect 331954 133378 331986 133614
rect 332222 133378 332306 133614
rect 332542 133378 332574 133614
rect 331954 133294 332574 133378
rect 331954 133058 331986 133294
rect 332222 133058 332306 133294
rect 332542 133058 332574 133294
rect 331954 93614 332574 133058
rect 331954 93378 331986 93614
rect 332222 93378 332306 93614
rect 332542 93378 332574 93614
rect 331954 93294 332574 93378
rect 331954 93058 331986 93294
rect 332222 93058 332306 93294
rect 332542 93058 332574 93294
rect 331954 53614 332574 93058
rect 331954 53378 331986 53614
rect 332222 53378 332306 53614
rect 332542 53378 332574 53614
rect 331954 53294 332574 53378
rect 331954 53058 331986 53294
rect 332222 53058 332306 53294
rect 332542 53058 332574 53294
rect 331954 13614 332574 53058
rect 331954 13378 331986 13614
rect 332222 13378 332306 13614
rect 332542 13378 332574 13614
rect 331954 13294 332574 13378
rect 331954 13058 331986 13294
rect 332222 13058 332306 13294
rect 332542 13058 332574 13294
rect 311954 -7302 311986 -7066
rect 312222 -7302 312306 -7066
rect 312542 -7302 312574 -7066
rect 311954 -7386 312574 -7302
rect 311954 -7622 311986 -7386
rect 312222 -7622 312306 -7386
rect 312542 -7622 312574 -7386
rect 311954 -7654 312574 -7622
rect 331954 -6106 332574 13058
rect 340794 705798 341414 705830
rect 340794 705562 340826 705798
rect 341062 705562 341146 705798
rect 341382 705562 341414 705798
rect 340794 705478 341414 705562
rect 340794 705242 340826 705478
rect 341062 705242 341146 705478
rect 341382 705242 341414 705478
rect 340794 662454 341414 705242
rect 340794 662218 340826 662454
rect 341062 662218 341146 662454
rect 341382 662218 341414 662454
rect 340794 662134 341414 662218
rect 340794 661898 340826 662134
rect 341062 661898 341146 662134
rect 341382 661898 341414 662134
rect 340794 622454 341414 661898
rect 340794 622218 340826 622454
rect 341062 622218 341146 622454
rect 341382 622218 341414 622454
rect 340794 622134 341414 622218
rect 340794 621898 340826 622134
rect 341062 621898 341146 622134
rect 341382 621898 341414 622134
rect 340794 582454 341414 621898
rect 340794 582218 340826 582454
rect 341062 582218 341146 582454
rect 341382 582218 341414 582454
rect 340794 582134 341414 582218
rect 340794 581898 340826 582134
rect 341062 581898 341146 582134
rect 341382 581898 341414 582134
rect 340794 542454 341414 581898
rect 340794 542218 340826 542454
rect 341062 542218 341146 542454
rect 341382 542218 341414 542454
rect 340794 542134 341414 542218
rect 340794 541898 340826 542134
rect 341062 541898 341146 542134
rect 341382 541898 341414 542134
rect 340794 502454 341414 541898
rect 340794 502218 340826 502454
rect 341062 502218 341146 502454
rect 341382 502218 341414 502454
rect 340794 502134 341414 502218
rect 340794 501898 340826 502134
rect 341062 501898 341146 502134
rect 341382 501898 341414 502134
rect 340794 462454 341414 501898
rect 340794 462218 340826 462454
rect 341062 462218 341146 462454
rect 341382 462218 341414 462454
rect 340794 462134 341414 462218
rect 340794 461898 340826 462134
rect 341062 461898 341146 462134
rect 341382 461898 341414 462134
rect 340794 422454 341414 461898
rect 340794 422218 340826 422454
rect 341062 422218 341146 422454
rect 341382 422218 341414 422454
rect 340794 422134 341414 422218
rect 340794 421898 340826 422134
rect 341062 421898 341146 422134
rect 341382 421898 341414 422134
rect 340794 382454 341414 421898
rect 340794 382218 340826 382454
rect 341062 382218 341146 382454
rect 341382 382218 341414 382454
rect 340794 382134 341414 382218
rect 340794 381898 340826 382134
rect 341062 381898 341146 382134
rect 341382 381898 341414 382134
rect 340794 342454 341414 381898
rect 340794 342218 340826 342454
rect 341062 342218 341146 342454
rect 341382 342218 341414 342454
rect 340794 342134 341414 342218
rect 340794 341898 340826 342134
rect 341062 341898 341146 342134
rect 341382 341898 341414 342134
rect 340794 302454 341414 341898
rect 340794 302218 340826 302454
rect 341062 302218 341146 302454
rect 341382 302218 341414 302454
rect 340794 302134 341414 302218
rect 340794 301898 340826 302134
rect 341062 301898 341146 302134
rect 341382 301898 341414 302134
rect 340794 262454 341414 301898
rect 340794 262218 340826 262454
rect 341062 262218 341146 262454
rect 341382 262218 341414 262454
rect 340794 262134 341414 262218
rect 340794 261898 340826 262134
rect 341062 261898 341146 262134
rect 341382 261898 341414 262134
rect 340794 222454 341414 261898
rect 340794 222218 340826 222454
rect 341062 222218 341146 222454
rect 341382 222218 341414 222454
rect 340794 222134 341414 222218
rect 340794 221898 340826 222134
rect 341062 221898 341146 222134
rect 341382 221898 341414 222134
rect 340794 182454 341414 221898
rect 340794 182218 340826 182454
rect 341062 182218 341146 182454
rect 341382 182218 341414 182454
rect 340794 182134 341414 182218
rect 340794 181898 340826 182134
rect 341062 181898 341146 182134
rect 341382 181898 341414 182134
rect 340794 142454 341414 181898
rect 340794 142218 340826 142454
rect 341062 142218 341146 142454
rect 341382 142218 341414 142454
rect 340794 142134 341414 142218
rect 340794 141898 340826 142134
rect 341062 141898 341146 142134
rect 341382 141898 341414 142134
rect 340794 102454 341414 141898
rect 340794 102218 340826 102454
rect 341062 102218 341146 102454
rect 341382 102218 341414 102454
rect 340794 102134 341414 102218
rect 340794 101898 340826 102134
rect 341062 101898 341146 102134
rect 341382 101898 341414 102134
rect 340794 62454 341414 101898
rect 340794 62218 340826 62454
rect 341062 62218 341146 62454
rect 341382 62218 341414 62454
rect 340794 62134 341414 62218
rect 340794 61898 340826 62134
rect 341062 61898 341146 62134
rect 341382 61898 341414 62134
rect 340794 22454 341414 61898
rect 340794 22218 340826 22454
rect 341062 22218 341146 22454
rect 341382 22218 341414 22454
rect 340794 22134 341414 22218
rect 340794 21898 340826 22134
rect 341062 21898 341146 22134
rect 341382 21898 341414 22134
rect 340794 -1306 341414 21898
rect 340794 -1542 340826 -1306
rect 341062 -1542 341146 -1306
rect 341382 -1542 341414 -1306
rect 340794 -1626 341414 -1542
rect 340794 -1862 340826 -1626
rect 341062 -1862 341146 -1626
rect 341382 -1862 341414 -1626
rect 340794 -1894 341414 -1862
rect 344514 666174 345134 707162
rect 344514 665938 344546 666174
rect 344782 665938 344866 666174
rect 345102 665938 345134 666174
rect 344514 665854 345134 665938
rect 344514 665618 344546 665854
rect 344782 665618 344866 665854
rect 345102 665618 345134 665854
rect 344514 626174 345134 665618
rect 344514 625938 344546 626174
rect 344782 625938 344866 626174
rect 345102 625938 345134 626174
rect 344514 625854 345134 625938
rect 344514 625618 344546 625854
rect 344782 625618 344866 625854
rect 345102 625618 345134 625854
rect 344514 586174 345134 625618
rect 344514 585938 344546 586174
rect 344782 585938 344866 586174
rect 345102 585938 345134 586174
rect 344514 585854 345134 585938
rect 344514 585618 344546 585854
rect 344782 585618 344866 585854
rect 345102 585618 345134 585854
rect 344514 546174 345134 585618
rect 344514 545938 344546 546174
rect 344782 545938 344866 546174
rect 345102 545938 345134 546174
rect 344514 545854 345134 545938
rect 344514 545618 344546 545854
rect 344782 545618 344866 545854
rect 345102 545618 345134 545854
rect 344514 506174 345134 545618
rect 344514 505938 344546 506174
rect 344782 505938 344866 506174
rect 345102 505938 345134 506174
rect 344514 505854 345134 505938
rect 344514 505618 344546 505854
rect 344782 505618 344866 505854
rect 345102 505618 345134 505854
rect 344514 466174 345134 505618
rect 344514 465938 344546 466174
rect 344782 465938 344866 466174
rect 345102 465938 345134 466174
rect 344514 465854 345134 465938
rect 344514 465618 344546 465854
rect 344782 465618 344866 465854
rect 345102 465618 345134 465854
rect 344514 426174 345134 465618
rect 344514 425938 344546 426174
rect 344782 425938 344866 426174
rect 345102 425938 345134 426174
rect 344514 425854 345134 425938
rect 344514 425618 344546 425854
rect 344782 425618 344866 425854
rect 345102 425618 345134 425854
rect 344514 386174 345134 425618
rect 344514 385938 344546 386174
rect 344782 385938 344866 386174
rect 345102 385938 345134 386174
rect 344514 385854 345134 385938
rect 344514 385618 344546 385854
rect 344782 385618 344866 385854
rect 345102 385618 345134 385854
rect 344514 346174 345134 385618
rect 344514 345938 344546 346174
rect 344782 345938 344866 346174
rect 345102 345938 345134 346174
rect 344514 345854 345134 345938
rect 344514 345618 344546 345854
rect 344782 345618 344866 345854
rect 345102 345618 345134 345854
rect 344514 306174 345134 345618
rect 344514 305938 344546 306174
rect 344782 305938 344866 306174
rect 345102 305938 345134 306174
rect 344514 305854 345134 305938
rect 344514 305618 344546 305854
rect 344782 305618 344866 305854
rect 345102 305618 345134 305854
rect 344514 266174 345134 305618
rect 344514 265938 344546 266174
rect 344782 265938 344866 266174
rect 345102 265938 345134 266174
rect 344514 265854 345134 265938
rect 344514 265618 344546 265854
rect 344782 265618 344866 265854
rect 345102 265618 345134 265854
rect 344514 226174 345134 265618
rect 344514 225938 344546 226174
rect 344782 225938 344866 226174
rect 345102 225938 345134 226174
rect 344514 225854 345134 225938
rect 344514 225618 344546 225854
rect 344782 225618 344866 225854
rect 345102 225618 345134 225854
rect 344514 186174 345134 225618
rect 344514 185938 344546 186174
rect 344782 185938 344866 186174
rect 345102 185938 345134 186174
rect 344514 185854 345134 185938
rect 344514 185618 344546 185854
rect 344782 185618 344866 185854
rect 345102 185618 345134 185854
rect 344514 146174 345134 185618
rect 344514 145938 344546 146174
rect 344782 145938 344866 146174
rect 345102 145938 345134 146174
rect 344514 145854 345134 145938
rect 344514 145618 344546 145854
rect 344782 145618 344866 145854
rect 345102 145618 345134 145854
rect 344514 106174 345134 145618
rect 344514 105938 344546 106174
rect 344782 105938 344866 106174
rect 345102 105938 345134 106174
rect 344514 105854 345134 105938
rect 344514 105618 344546 105854
rect 344782 105618 344866 105854
rect 345102 105618 345134 105854
rect 344514 66174 345134 105618
rect 344514 65938 344546 66174
rect 344782 65938 344866 66174
rect 345102 65938 345134 66174
rect 344514 65854 345134 65938
rect 344514 65618 344546 65854
rect 344782 65618 344866 65854
rect 345102 65618 345134 65854
rect 344514 26174 345134 65618
rect 344514 25938 344546 26174
rect 344782 25938 344866 26174
rect 345102 25938 345134 26174
rect 344514 25854 345134 25938
rect 344514 25618 344546 25854
rect 344782 25618 344866 25854
rect 345102 25618 345134 25854
rect 344514 -3226 345134 25618
rect 344514 -3462 344546 -3226
rect 344782 -3462 344866 -3226
rect 345102 -3462 345134 -3226
rect 344514 -3546 345134 -3462
rect 344514 -3782 344546 -3546
rect 344782 -3782 344866 -3546
rect 345102 -3782 345134 -3546
rect 344514 -3814 345134 -3782
rect 348234 669894 348854 709082
rect 348234 669658 348266 669894
rect 348502 669658 348586 669894
rect 348822 669658 348854 669894
rect 348234 669574 348854 669658
rect 348234 669338 348266 669574
rect 348502 669338 348586 669574
rect 348822 669338 348854 669574
rect 348234 629894 348854 669338
rect 348234 629658 348266 629894
rect 348502 629658 348586 629894
rect 348822 629658 348854 629894
rect 348234 629574 348854 629658
rect 348234 629338 348266 629574
rect 348502 629338 348586 629574
rect 348822 629338 348854 629574
rect 348234 589894 348854 629338
rect 348234 589658 348266 589894
rect 348502 589658 348586 589894
rect 348822 589658 348854 589894
rect 348234 589574 348854 589658
rect 348234 589338 348266 589574
rect 348502 589338 348586 589574
rect 348822 589338 348854 589574
rect 348234 549894 348854 589338
rect 348234 549658 348266 549894
rect 348502 549658 348586 549894
rect 348822 549658 348854 549894
rect 348234 549574 348854 549658
rect 348234 549338 348266 549574
rect 348502 549338 348586 549574
rect 348822 549338 348854 549574
rect 348234 509894 348854 549338
rect 348234 509658 348266 509894
rect 348502 509658 348586 509894
rect 348822 509658 348854 509894
rect 348234 509574 348854 509658
rect 348234 509338 348266 509574
rect 348502 509338 348586 509574
rect 348822 509338 348854 509574
rect 348234 469894 348854 509338
rect 348234 469658 348266 469894
rect 348502 469658 348586 469894
rect 348822 469658 348854 469894
rect 348234 469574 348854 469658
rect 348234 469338 348266 469574
rect 348502 469338 348586 469574
rect 348822 469338 348854 469574
rect 348234 429894 348854 469338
rect 348234 429658 348266 429894
rect 348502 429658 348586 429894
rect 348822 429658 348854 429894
rect 348234 429574 348854 429658
rect 348234 429338 348266 429574
rect 348502 429338 348586 429574
rect 348822 429338 348854 429574
rect 348234 389894 348854 429338
rect 348234 389658 348266 389894
rect 348502 389658 348586 389894
rect 348822 389658 348854 389894
rect 348234 389574 348854 389658
rect 348234 389338 348266 389574
rect 348502 389338 348586 389574
rect 348822 389338 348854 389574
rect 348234 349894 348854 389338
rect 348234 349658 348266 349894
rect 348502 349658 348586 349894
rect 348822 349658 348854 349894
rect 348234 349574 348854 349658
rect 348234 349338 348266 349574
rect 348502 349338 348586 349574
rect 348822 349338 348854 349574
rect 348234 309894 348854 349338
rect 348234 309658 348266 309894
rect 348502 309658 348586 309894
rect 348822 309658 348854 309894
rect 348234 309574 348854 309658
rect 348234 309338 348266 309574
rect 348502 309338 348586 309574
rect 348822 309338 348854 309574
rect 348234 269894 348854 309338
rect 348234 269658 348266 269894
rect 348502 269658 348586 269894
rect 348822 269658 348854 269894
rect 348234 269574 348854 269658
rect 348234 269338 348266 269574
rect 348502 269338 348586 269574
rect 348822 269338 348854 269574
rect 348234 229894 348854 269338
rect 348234 229658 348266 229894
rect 348502 229658 348586 229894
rect 348822 229658 348854 229894
rect 348234 229574 348854 229658
rect 348234 229338 348266 229574
rect 348502 229338 348586 229574
rect 348822 229338 348854 229574
rect 348234 189894 348854 229338
rect 348234 189658 348266 189894
rect 348502 189658 348586 189894
rect 348822 189658 348854 189894
rect 348234 189574 348854 189658
rect 348234 189338 348266 189574
rect 348502 189338 348586 189574
rect 348822 189338 348854 189574
rect 348234 149894 348854 189338
rect 348234 149658 348266 149894
rect 348502 149658 348586 149894
rect 348822 149658 348854 149894
rect 348234 149574 348854 149658
rect 348234 149338 348266 149574
rect 348502 149338 348586 149574
rect 348822 149338 348854 149574
rect 348234 109894 348854 149338
rect 348234 109658 348266 109894
rect 348502 109658 348586 109894
rect 348822 109658 348854 109894
rect 348234 109574 348854 109658
rect 348234 109338 348266 109574
rect 348502 109338 348586 109574
rect 348822 109338 348854 109574
rect 348234 69894 348854 109338
rect 348234 69658 348266 69894
rect 348502 69658 348586 69894
rect 348822 69658 348854 69894
rect 348234 69574 348854 69658
rect 348234 69338 348266 69574
rect 348502 69338 348586 69574
rect 348822 69338 348854 69574
rect 348234 29894 348854 69338
rect 348234 29658 348266 29894
rect 348502 29658 348586 29894
rect 348822 29658 348854 29894
rect 348234 29574 348854 29658
rect 348234 29338 348266 29574
rect 348502 29338 348586 29574
rect 348822 29338 348854 29574
rect 348234 -5146 348854 29338
rect 348234 -5382 348266 -5146
rect 348502 -5382 348586 -5146
rect 348822 -5382 348854 -5146
rect 348234 -5466 348854 -5382
rect 348234 -5702 348266 -5466
rect 348502 -5702 348586 -5466
rect 348822 -5702 348854 -5466
rect 348234 -5734 348854 -5702
rect 351954 673614 352574 711002
rect 371954 710598 372574 711590
rect 371954 710362 371986 710598
rect 372222 710362 372306 710598
rect 372542 710362 372574 710598
rect 371954 710278 372574 710362
rect 371954 710042 371986 710278
rect 372222 710042 372306 710278
rect 372542 710042 372574 710278
rect 368234 708678 368854 709670
rect 368234 708442 368266 708678
rect 368502 708442 368586 708678
rect 368822 708442 368854 708678
rect 368234 708358 368854 708442
rect 368234 708122 368266 708358
rect 368502 708122 368586 708358
rect 368822 708122 368854 708358
rect 364514 706758 365134 707750
rect 364514 706522 364546 706758
rect 364782 706522 364866 706758
rect 365102 706522 365134 706758
rect 364514 706438 365134 706522
rect 364514 706202 364546 706438
rect 364782 706202 364866 706438
rect 365102 706202 365134 706438
rect 351954 673378 351986 673614
rect 352222 673378 352306 673614
rect 352542 673378 352574 673614
rect 351954 673294 352574 673378
rect 351954 673058 351986 673294
rect 352222 673058 352306 673294
rect 352542 673058 352574 673294
rect 351954 633614 352574 673058
rect 351954 633378 351986 633614
rect 352222 633378 352306 633614
rect 352542 633378 352574 633614
rect 351954 633294 352574 633378
rect 351954 633058 351986 633294
rect 352222 633058 352306 633294
rect 352542 633058 352574 633294
rect 351954 593614 352574 633058
rect 351954 593378 351986 593614
rect 352222 593378 352306 593614
rect 352542 593378 352574 593614
rect 351954 593294 352574 593378
rect 351954 593058 351986 593294
rect 352222 593058 352306 593294
rect 352542 593058 352574 593294
rect 351954 553614 352574 593058
rect 351954 553378 351986 553614
rect 352222 553378 352306 553614
rect 352542 553378 352574 553614
rect 351954 553294 352574 553378
rect 351954 553058 351986 553294
rect 352222 553058 352306 553294
rect 352542 553058 352574 553294
rect 351954 513614 352574 553058
rect 351954 513378 351986 513614
rect 352222 513378 352306 513614
rect 352542 513378 352574 513614
rect 351954 513294 352574 513378
rect 351954 513058 351986 513294
rect 352222 513058 352306 513294
rect 352542 513058 352574 513294
rect 351954 473614 352574 513058
rect 351954 473378 351986 473614
rect 352222 473378 352306 473614
rect 352542 473378 352574 473614
rect 351954 473294 352574 473378
rect 351954 473058 351986 473294
rect 352222 473058 352306 473294
rect 352542 473058 352574 473294
rect 351954 433614 352574 473058
rect 351954 433378 351986 433614
rect 352222 433378 352306 433614
rect 352542 433378 352574 433614
rect 351954 433294 352574 433378
rect 351954 433058 351986 433294
rect 352222 433058 352306 433294
rect 352542 433058 352574 433294
rect 351954 393614 352574 433058
rect 351954 393378 351986 393614
rect 352222 393378 352306 393614
rect 352542 393378 352574 393614
rect 351954 393294 352574 393378
rect 351954 393058 351986 393294
rect 352222 393058 352306 393294
rect 352542 393058 352574 393294
rect 351954 353614 352574 393058
rect 351954 353378 351986 353614
rect 352222 353378 352306 353614
rect 352542 353378 352574 353614
rect 351954 353294 352574 353378
rect 351954 353058 351986 353294
rect 352222 353058 352306 353294
rect 352542 353058 352574 353294
rect 351954 313614 352574 353058
rect 351954 313378 351986 313614
rect 352222 313378 352306 313614
rect 352542 313378 352574 313614
rect 351954 313294 352574 313378
rect 351954 313058 351986 313294
rect 352222 313058 352306 313294
rect 352542 313058 352574 313294
rect 351954 273614 352574 313058
rect 351954 273378 351986 273614
rect 352222 273378 352306 273614
rect 352542 273378 352574 273614
rect 351954 273294 352574 273378
rect 351954 273058 351986 273294
rect 352222 273058 352306 273294
rect 352542 273058 352574 273294
rect 351954 233614 352574 273058
rect 351954 233378 351986 233614
rect 352222 233378 352306 233614
rect 352542 233378 352574 233614
rect 351954 233294 352574 233378
rect 351954 233058 351986 233294
rect 352222 233058 352306 233294
rect 352542 233058 352574 233294
rect 351954 193614 352574 233058
rect 351954 193378 351986 193614
rect 352222 193378 352306 193614
rect 352542 193378 352574 193614
rect 351954 193294 352574 193378
rect 351954 193058 351986 193294
rect 352222 193058 352306 193294
rect 352542 193058 352574 193294
rect 351954 153614 352574 193058
rect 351954 153378 351986 153614
rect 352222 153378 352306 153614
rect 352542 153378 352574 153614
rect 351954 153294 352574 153378
rect 351954 153058 351986 153294
rect 352222 153058 352306 153294
rect 352542 153058 352574 153294
rect 351954 113614 352574 153058
rect 351954 113378 351986 113614
rect 352222 113378 352306 113614
rect 352542 113378 352574 113614
rect 351954 113294 352574 113378
rect 351954 113058 351986 113294
rect 352222 113058 352306 113294
rect 352542 113058 352574 113294
rect 351954 73614 352574 113058
rect 351954 73378 351986 73614
rect 352222 73378 352306 73614
rect 352542 73378 352574 73614
rect 351954 73294 352574 73378
rect 351954 73058 351986 73294
rect 352222 73058 352306 73294
rect 352542 73058 352574 73294
rect 351954 33614 352574 73058
rect 351954 33378 351986 33614
rect 352222 33378 352306 33614
rect 352542 33378 352574 33614
rect 351954 33294 352574 33378
rect 351954 33058 351986 33294
rect 352222 33058 352306 33294
rect 352542 33058 352574 33294
rect 331954 -6342 331986 -6106
rect 332222 -6342 332306 -6106
rect 332542 -6342 332574 -6106
rect 331954 -6426 332574 -6342
rect 331954 -6662 331986 -6426
rect 332222 -6662 332306 -6426
rect 332542 -6662 332574 -6426
rect 331954 -7654 332574 -6662
rect 351954 -7066 352574 33058
rect 360794 704838 361414 705830
rect 360794 704602 360826 704838
rect 361062 704602 361146 704838
rect 361382 704602 361414 704838
rect 360794 704518 361414 704602
rect 360794 704282 360826 704518
rect 361062 704282 361146 704518
rect 361382 704282 361414 704518
rect 360794 682454 361414 704282
rect 360794 682218 360826 682454
rect 361062 682218 361146 682454
rect 361382 682218 361414 682454
rect 360794 682134 361414 682218
rect 360794 681898 360826 682134
rect 361062 681898 361146 682134
rect 361382 681898 361414 682134
rect 360794 642454 361414 681898
rect 360794 642218 360826 642454
rect 361062 642218 361146 642454
rect 361382 642218 361414 642454
rect 360794 642134 361414 642218
rect 360794 641898 360826 642134
rect 361062 641898 361146 642134
rect 361382 641898 361414 642134
rect 360794 602454 361414 641898
rect 360794 602218 360826 602454
rect 361062 602218 361146 602454
rect 361382 602218 361414 602454
rect 360794 602134 361414 602218
rect 360794 601898 360826 602134
rect 361062 601898 361146 602134
rect 361382 601898 361414 602134
rect 360794 562454 361414 601898
rect 360794 562218 360826 562454
rect 361062 562218 361146 562454
rect 361382 562218 361414 562454
rect 360794 562134 361414 562218
rect 360794 561898 360826 562134
rect 361062 561898 361146 562134
rect 361382 561898 361414 562134
rect 360794 522454 361414 561898
rect 360794 522218 360826 522454
rect 361062 522218 361146 522454
rect 361382 522218 361414 522454
rect 360794 522134 361414 522218
rect 360794 521898 360826 522134
rect 361062 521898 361146 522134
rect 361382 521898 361414 522134
rect 360794 482454 361414 521898
rect 360794 482218 360826 482454
rect 361062 482218 361146 482454
rect 361382 482218 361414 482454
rect 360794 482134 361414 482218
rect 360794 481898 360826 482134
rect 361062 481898 361146 482134
rect 361382 481898 361414 482134
rect 360794 442454 361414 481898
rect 360794 442218 360826 442454
rect 361062 442218 361146 442454
rect 361382 442218 361414 442454
rect 360794 442134 361414 442218
rect 360794 441898 360826 442134
rect 361062 441898 361146 442134
rect 361382 441898 361414 442134
rect 360794 402454 361414 441898
rect 360794 402218 360826 402454
rect 361062 402218 361146 402454
rect 361382 402218 361414 402454
rect 360794 402134 361414 402218
rect 360794 401898 360826 402134
rect 361062 401898 361146 402134
rect 361382 401898 361414 402134
rect 360794 362454 361414 401898
rect 360794 362218 360826 362454
rect 361062 362218 361146 362454
rect 361382 362218 361414 362454
rect 360794 362134 361414 362218
rect 360794 361898 360826 362134
rect 361062 361898 361146 362134
rect 361382 361898 361414 362134
rect 360794 322454 361414 361898
rect 360794 322218 360826 322454
rect 361062 322218 361146 322454
rect 361382 322218 361414 322454
rect 360794 322134 361414 322218
rect 360794 321898 360826 322134
rect 361062 321898 361146 322134
rect 361382 321898 361414 322134
rect 360794 282454 361414 321898
rect 360794 282218 360826 282454
rect 361062 282218 361146 282454
rect 361382 282218 361414 282454
rect 360794 282134 361414 282218
rect 360794 281898 360826 282134
rect 361062 281898 361146 282134
rect 361382 281898 361414 282134
rect 360794 242454 361414 281898
rect 360794 242218 360826 242454
rect 361062 242218 361146 242454
rect 361382 242218 361414 242454
rect 360794 242134 361414 242218
rect 360794 241898 360826 242134
rect 361062 241898 361146 242134
rect 361382 241898 361414 242134
rect 360794 202454 361414 241898
rect 360794 202218 360826 202454
rect 361062 202218 361146 202454
rect 361382 202218 361414 202454
rect 360794 202134 361414 202218
rect 360794 201898 360826 202134
rect 361062 201898 361146 202134
rect 361382 201898 361414 202134
rect 360794 162454 361414 201898
rect 360794 162218 360826 162454
rect 361062 162218 361146 162454
rect 361382 162218 361414 162454
rect 360794 162134 361414 162218
rect 360794 161898 360826 162134
rect 361062 161898 361146 162134
rect 361382 161898 361414 162134
rect 360794 122454 361414 161898
rect 360794 122218 360826 122454
rect 361062 122218 361146 122454
rect 361382 122218 361414 122454
rect 360794 122134 361414 122218
rect 360794 121898 360826 122134
rect 361062 121898 361146 122134
rect 361382 121898 361414 122134
rect 360794 82454 361414 121898
rect 360794 82218 360826 82454
rect 361062 82218 361146 82454
rect 361382 82218 361414 82454
rect 360794 82134 361414 82218
rect 360794 81898 360826 82134
rect 361062 81898 361146 82134
rect 361382 81898 361414 82134
rect 360794 42454 361414 81898
rect 360794 42218 360826 42454
rect 361062 42218 361146 42454
rect 361382 42218 361414 42454
rect 360794 42134 361414 42218
rect 360794 41898 360826 42134
rect 361062 41898 361146 42134
rect 361382 41898 361414 42134
rect 360794 2454 361414 41898
rect 360794 2218 360826 2454
rect 361062 2218 361146 2454
rect 361382 2218 361414 2454
rect 360794 2134 361414 2218
rect 360794 1898 360826 2134
rect 361062 1898 361146 2134
rect 361382 1898 361414 2134
rect 360794 -346 361414 1898
rect 360794 -582 360826 -346
rect 361062 -582 361146 -346
rect 361382 -582 361414 -346
rect 360794 -666 361414 -582
rect 360794 -902 360826 -666
rect 361062 -902 361146 -666
rect 361382 -902 361414 -666
rect 360794 -1894 361414 -902
rect 364514 686174 365134 706202
rect 364514 685938 364546 686174
rect 364782 685938 364866 686174
rect 365102 685938 365134 686174
rect 364514 685854 365134 685938
rect 364514 685618 364546 685854
rect 364782 685618 364866 685854
rect 365102 685618 365134 685854
rect 364514 646174 365134 685618
rect 364514 645938 364546 646174
rect 364782 645938 364866 646174
rect 365102 645938 365134 646174
rect 364514 645854 365134 645938
rect 364514 645618 364546 645854
rect 364782 645618 364866 645854
rect 365102 645618 365134 645854
rect 364514 606174 365134 645618
rect 364514 605938 364546 606174
rect 364782 605938 364866 606174
rect 365102 605938 365134 606174
rect 364514 605854 365134 605938
rect 364514 605618 364546 605854
rect 364782 605618 364866 605854
rect 365102 605618 365134 605854
rect 364514 566174 365134 605618
rect 364514 565938 364546 566174
rect 364782 565938 364866 566174
rect 365102 565938 365134 566174
rect 364514 565854 365134 565938
rect 364514 565618 364546 565854
rect 364782 565618 364866 565854
rect 365102 565618 365134 565854
rect 364514 526174 365134 565618
rect 364514 525938 364546 526174
rect 364782 525938 364866 526174
rect 365102 525938 365134 526174
rect 364514 525854 365134 525938
rect 364514 525618 364546 525854
rect 364782 525618 364866 525854
rect 365102 525618 365134 525854
rect 364514 486174 365134 525618
rect 364514 485938 364546 486174
rect 364782 485938 364866 486174
rect 365102 485938 365134 486174
rect 364514 485854 365134 485938
rect 364514 485618 364546 485854
rect 364782 485618 364866 485854
rect 365102 485618 365134 485854
rect 364514 446174 365134 485618
rect 364514 445938 364546 446174
rect 364782 445938 364866 446174
rect 365102 445938 365134 446174
rect 364514 445854 365134 445938
rect 364514 445618 364546 445854
rect 364782 445618 364866 445854
rect 365102 445618 365134 445854
rect 364514 406174 365134 445618
rect 364514 405938 364546 406174
rect 364782 405938 364866 406174
rect 365102 405938 365134 406174
rect 364514 405854 365134 405938
rect 364514 405618 364546 405854
rect 364782 405618 364866 405854
rect 365102 405618 365134 405854
rect 364514 366174 365134 405618
rect 364514 365938 364546 366174
rect 364782 365938 364866 366174
rect 365102 365938 365134 366174
rect 364514 365854 365134 365938
rect 364514 365618 364546 365854
rect 364782 365618 364866 365854
rect 365102 365618 365134 365854
rect 364514 326174 365134 365618
rect 364514 325938 364546 326174
rect 364782 325938 364866 326174
rect 365102 325938 365134 326174
rect 364514 325854 365134 325938
rect 364514 325618 364546 325854
rect 364782 325618 364866 325854
rect 365102 325618 365134 325854
rect 364514 286174 365134 325618
rect 364514 285938 364546 286174
rect 364782 285938 364866 286174
rect 365102 285938 365134 286174
rect 364514 285854 365134 285938
rect 364514 285618 364546 285854
rect 364782 285618 364866 285854
rect 365102 285618 365134 285854
rect 364514 246174 365134 285618
rect 364514 245938 364546 246174
rect 364782 245938 364866 246174
rect 365102 245938 365134 246174
rect 364514 245854 365134 245938
rect 364514 245618 364546 245854
rect 364782 245618 364866 245854
rect 365102 245618 365134 245854
rect 364514 206174 365134 245618
rect 364514 205938 364546 206174
rect 364782 205938 364866 206174
rect 365102 205938 365134 206174
rect 364514 205854 365134 205938
rect 364514 205618 364546 205854
rect 364782 205618 364866 205854
rect 365102 205618 365134 205854
rect 364514 166174 365134 205618
rect 364514 165938 364546 166174
rect 364782 165938 364866 166174
rect 365102 165938 365134 166174
rect 364514 165854 365134 165938
rect 364514 165618 364546 165854
rect 364782 165618 364866 165854
rect 365102 165618 365134 165854
rect 364514 126174 365134 165618
rect 364514 125938 364546 126174
rect 364782 125938 364866 126174
rect 365102 125938 365134 126174
rect 364514 125854 365134 125938
rect 364514 125618 364546 125854
rect 364782 125618 364866 125854
rect 365102 125618 365134 125854
rect 364514 86174 365134 125618
rect 364514 85938 364546 86174
rect 364782 85938 364866 86174
rect 365102 85938 365134 86174
rect 364514 85854 365134 85938
rect 364514 85618 364546 85854
rect 364782 85618 364866 85854
rect 365102 85618 365134 85854
rect 364514 46174 365134 85618
rect 364514 45938 364546 46174
rect 364782 45938 364866 46174
rect 365102 45938 365134 46174
rect 364514 45854 365134 45938
rect 364514 45618 364546 45854
rect 364782 45618 364866 45854
rect 365102 45618 365134 45854
rect 364514 6174 365134 45618
rect 364514 5938 364546 6174
rect 364782 5938 364866 6174
rect 365102 5938 365134 6174
rect 364514 5854 365134 5938
rect 364514 5618 364546 5854
rect 364782 5618 364866 5854
rect 365102 5618 365134 5854
rect 364514 -2266 365134 5618
rect 364514 -2502 364546 -2266
rect 364782 -2502 364866 -2266
rect 365102 -2502 365134 -2266
rect 364514 -2586 365134 -2502
rect 364514 -2822 364546 -2586
rect 364782 -2822 364866 -2586
rect 365102 -2822 365134 -2586
rect 364514 -3814 365134 -2822
rect 368234 689894 368854 708122
rect 368234 689658 368266 689894
rect 368502 689658 368586 689894
rect 368822 689658 368854 689894
rect 368234 689574 368854 689658
rect 368234 689338 368266 689574
rect 368502 689338 368586 689574
rect 368822 689338 368854 689574
rect 368234 649894 368854 689338
rect 368234 649658 368266 649894
rect 368502 649658 368586 649894
rect 368822 649658 368854 649894
rect 368234 649574 368854 649658
rect 368234 649338 368266 649574
rect 368502 649338 368586 649574
rect 368822 649338 368854 649574
rect 368234 609894 368854 649338
rect 368234 609658 368266 609894
rect 368502 609658 368586 609894
rect 368822 609658 368854 609894
rect 368234 609574 368854 609658
rect 368234 609338 368266 609574
rect 368502 609338 368586 609574
rect 368822 609338 368854 609574
rect 368234 569894 368854 609338
rect 368234 569658 368266 569894
rect 368502 569658 368586 569894
rect 368822 569658 368854 569894
rect 368234 569574 368854 569658
rect 368234 569338 368266 569574
rect 368502 569338 368586 569574
rect 368822 569338 368854 569574
rect 368234 529894 368854 569338
rect 368234 529658 368266 529894
rect 368502 529658 368586 529894
rect 368822 529658 368854 529894
rect 368234 529574 368854 529658
rect 368234 529338 368266 529574
rect 368502 529338 368586 529574
rect 368822 529338 368854 529574
rect 368234 489894 368854 529338
rect 368234 489658 368266 489894
rect 368502 489658 368586 489894
rect 368822 489658 368854 489894
rect 368234 489574 368854 489658
rect 368234 489338 368266 489574
rect 368502 489338 368586 489574
rect 368822 489338 368854 489574
rect 368234 449894 368854 489338
rect 368234 449658 368266 449894
rect 368502 449658 368586 449894
rect 368822 449658 368854 449894
rect 368234 449574 368854 449658
rect 368234 449338 368266 449574
rect 368502 449338 368586 449574
rect 368822 449338 368854 449574
rect 368234 409894 368854 449338
rect 368234 409658 368266 409894
rect 368502 409658 368586 409894
rect 368822 409658 368854 409894
rect 368234 409574 368854 409658
rect 368234 409338 368266 409574
rect 368502 409338 368586 409574
rect 368822 409338 368854 409574
rect 368234 369894 368854 409338
rect 368234 369658 368266 369894
rect 368502 369658 368586 369894
rect 368822 369658 368854 369894
rect 368234 369574 368854 369658
rect 368234 369338 368266 369574
rect 368502 369338 368586 369574
rect 368822 369338 368854 369574
rect 368234 329894 368854 369338
rect 368234 329658 368266 329894
rect 368502 329658 368586 329894
rect 368822 329658 368854 329894
rect 368234 329574 368854 329658
rect 368234 329338 368266 329574
rect 368502 329338 368586 329574
rect 368822 329338 368854 329574
rect 368234 289894 368854 329338
rect 368234 289658 368266 289894
rect 368502 289658 368586 289894
rect 368822 289658 368854 289894
rect 368234 289574 368854 289658
rect 368234 289338 368266 289574
rect 368502 289338 368586 289574
rect 368822 289338 368854 289574
rect 368234 249894 368854 289338
rect 368234 249658 368266 249894
rect 368502 249658 368586 249894
rect 368822 249658 368854 249894
rect 368234 249574 368854 249658
rect 368234 249338 368266 249574
rect 368502 249338 368586 249574
rect 368822 249338 368854 249574
rect 368234 209894 368854 249338
rect 368234 209658 368266 209894
rect 368502 209658 368586 209894
rect 368822 209658 368854 209894
rect 368234 209574 368854 209658
rect 368234 209338 368266 209574
rect 368502 209338 368586 209574
rect 368822 209338 368854 209574
rect 368234 169894 368854 209338
rect 368234 169658 368266 169894
rect 368502 169658 368586 169894
rect 368822 169658 368854 169894
rect 368234 169574 368854 169658
rect 368234 169338 368266 169574
rect 368502 169338 368586 169574
rect 368822 169338 368854 169574
rect 368234 129894 368854 169338
rect 368234 129658 368266 129894
rect 368502 129658 368586 129894
rect 368822 129658 368854 129894
rect 368234 129574 368854 129658
rect 368234 129338 368266 129574
rect 368502 129338 368586 129574
rect 368822 129338 368854 129574
rect 368234 89894 368854 129338
rect 368234 89658 368266 89894
rect 368502 89658 368586 89894
rect 368822 89658 368854 89894
rect 368234 89574 368854 89658
rect 368234 89338 368266 89574
rect 368502 89338 368586 89574
rect 368822 89338 368854 89574
rect 368234 49894 368854 89338
rect 368234 49658 368266 49894
rect 368502 49658 368586 49894
rect 368822 49658 368854 49894
rect 368234 49574 368854 49658
rect 368234 49338 368266 49574
rect 368502 49338 368586 49574
rect 368822 49338 368854 49574
rect 368234 9894 368854 49338
rect 368234 9658 368266 9894
rect 368502 9658 368586 9894
rect 368822 9658 368854 9894
rect 368234 9574 368854 9658
rect 368234 9338 368266 9574
rect 368502 9338 368586 9574
rect 368822 9338 368854 9574
rect 368234 -4186 368854 9338
rect 368234 -4422 368266 -4186
rect 368502 -4422 368586 -4186
rect 368822 -4422 368854 -4186
rect 368234 -4506 368854 -4422
rect 368234 -4742 368266 -4506
rect 368502 -4742 368586 -4506
rect 368822 -4742 368854 -4506
rect 368234 -5734 368854 -4742
rect 371954 693614 372574 710042
rect 391954 711558 392574 711590
rect 391954 711322 391986 711558
rect 392222 711322 392306 711558
rect 392542 711322 392574 711558
rect 391954 711238 392574 711322
rect 391954 711002 391986 711238
rect 392222 711002 392306 711238
rect 392542 711002 392574 711238
rect 388234 709638 388854 709670
rect 388234 709402 388266 709638
rect 388502 709402 388586 709638
rect 388822 709402 388854 709638
rect 388234 709318 388854 709402
rect 388234 709082 388266 709318
rect 388502 709082 388586 709318
rect 388822 709082 388854 709318
rect 384514 707718 385134 707750
rect 384514 707482 384546 707718
rect 384782 707482 384866 707718
rect 385102 707482 385134 707718
rect 384514 707398 385134 707482
rect 384514 707162 384546 707398
rect 384782 707162 384866 707398
rect 385102 707162 385134 707398
rect 371954 693378 371986 693614
rect 372222 693378 372306 693614
rect 372542 693378 372574 693614
rect 371954 693294 372574 693378
rect 371954 693058 371986 693294
rect 372222 693058 372306 693294
rect 372542 693058 372574 693294
rect 371954 653614 372574 693058
rect 371954 653378 371986 653614
rect 372222 653378 372306 653614
rect 372542 653378 372574 653614
rect 371954 653294 372574 653378
rect 371954 653058 371986 653294
rect 372222 653058 372306 653294
rect 372542 653058 372574 653294
rect 371954 613614 372574 653058
rect 371954 613378 371986 613614
rect 372222 613378 372306 613614
rect 372542 613378 372574 613614
rect 371954 613294 372574 613378
rect 371954 613058 371986 613294
rect 372222 613058 372306 613294
rect 372542 613058 372574 613294
rect 371954 573614 372574 613058
rect 371954 573378 371986 573614
rect 372222 573378 372306 573614
rect 372542 573378 372574 573614
rect 371954 573294 372574 573378
rect 371954 573058 371986 573294
rect 372222 573058 372306 573294
rect 372542 573058 372574 573294
rect 371954 533614 372574 573058
rect 371954 533378 371986 533614
rect 372222 533378 372306 533614
rect 372542 533378 372574 533614
rect 371954 533294 372574 533378
rect 371954 533058 371986 533294
rect 372222 533058 372306 533294
rect 372542 533058 372574 533294
rect 371954 493614 372574 533058
rect 371954 493378 371986 493614
rect 372222 493378 372306 493614
rect 372542 493378 372574 493614
rect 371954 493294 372574 493378
rect 371954 493058 371986 493294
rect 372222 493058 372306 493294
rect 372542 493058 372574 493294
rect 371954 453614 372574 493058
rect 371954 453378 371986 453614
rect 372222 453378 372306 453614
rect 372542 453378 372574 453614
rect 371954 453294 372574 453378
rect 371954 453058 371986 453294
rect 372222 453058 372306 453294
rect 372542 453058 372574 453294
rect 371954 413614 372574 453058
rect 371954 413378 371986 413614
rect 372222 413378 372306 413614
rect 372542 413378 372574 413614
rect 371954 413294 372574 413378
rect 371954 413058 371986 413294
rect 372222 413058 372306 413294
rect 372542 413058 372574 413294
rect 371954 373614 372574 413058
rect 371954 373378 371986 373614
rect 372222 373378 372306 373614
rect 372542 373378 372574 373614
rect 371954 373294 372574 373378
rect 371954 373058 371986 373294
rect 372222 373058 372306 373294
rect 372542 373058 372574 373294
rect 371954 333614 372574 373058
rect 371954 333378 371986 333614
rect 372222 333378 372306 333614
rect 372542 333378 372574 333614
rect 371954 333294 372574 333378
rect 371954 333058 371986 333294
rect 372222 333058 372306 333294
rect 372542 333058 372574 333294
rect 371954 293614 372574 333058
rect 371954 293378 371986 293614
rect 372222 293378 372306 293614
rect 372542 293378 372574 293614
rect 371954 293294 372574 293378
rect 371954 293058 371986 293294
rect 372222 293058 372306 293294
rect 372542 293058 372574 293294
rect 371954 253614 372574 293058
rect 371954 253378 371986 253614
rect 372222 253378 372306 253614
rect 372542 253378 372574 253614
rect 371954 253294 372574 253378
rect 371954 253058 371986 253294
rect 372222 253058 372306 253294
rect 372542 253058 372574 253294
rect 371954 213614 372574 253058
rect 371954 213378 371986 213614
rect 372222 213378 372306 213614
rect 372542 213378 372574 213614
rect 371954 213294 372574 213378
rect 371954 213058 371986 213294
rect 372222 213058 372306 213294
rect 372542 213058 372574 213294
rect 371954 173614 372574 213058
rect 371954 173378 371986 173614
rect 372222 173378 372306 173614
rect 372542 173378 372574 173614
rect 371954 173294 372574 173378
rect 371954 173058 371986 173294
rect 372222 173058 372306 173294
rect 372542 173058 372574 173294
rect 371954 133614 372574 173058
rect 371954 133378 371986 133614
rect 372222 133378 372306 133614
rect 372542 133378 372574 133614
rect 371954 133294 372574 133378
rect 371954 133058 371986 133294
rect 372222 133058 372306 133294
rect 372542 133058 372574 133294
rect 371954 93614 372574 133058
rect 371954 93378 371986 93614
rect 372222 93378 372306 93614
rect 372542 93378 372574 93614
rect 371954 93294 372574 93378
rect 371954 93058 371986 93294
rect 372222 93058 372306 93294
rect 372542 93058 372574 93294
rect 371954 53614 372574 93058
rect 371954 53378 371986 53614
rect 372222 53378 372306 53614
rect 372542 53378 372574 53614
rect 371954 53294 372574 53378
rect 371954 53058 371986 53294
rect 372222 53058 372306 53294
rect 372542 53058 372574 53294
rect 371954 13614 372574 53058
rect 371954 13378 371986 13614
rect 372222 13378 372306 13614
rect 372542 13378 372574 13614
rect 371954 13294 372574 13378
rect 371954 13058 371986 13294
rect 372222 13058 372306 13294
rect 372542 13058 372574 13294
rect 351954 -7302 351986 -7066
rect 352222 -7302 352306 -7066
rect 352542 -7302 352574 -7066
rect 351954 -7386 352574 -7302
rect 351954 -7622 351986 -7386
rect 352222 -7622 352306 -7386
rect 352542 -7622 352574 -7386
rect 351954 -7654 352574 -7622
rect 371954 -6106 372574 13058
rect 380794 705798 381414 705830
rect 380794 705562 380826 705798
rect 381062 705562 381146 705798
rect 381382 705562 381414 705798
rect 380794 705478 381414 705562
rect 380794 705242 380826 705478
rect 381062 705242 381146 705478
rect 381382 705242 381414 705478
rect 380794 662454 381414 705242
rect 380794 662218 380826 662454
rect 381062 662218 381146 662454
rect 381382 662218 381414 662454
rect 380794 662134 381414 662218
rect 380794 661898 380826 662134
rect 381062 661898 381146 662134
rect 381382 661898 381414 662134
rect 380794 622454 381414 661898
rect 380794 622218 380826 622454
rect 381062 622218 381146 622454
rect 381382 622218 381414 622454
rect 380794 622134 381414 622218
rect 380794 621898 380826 622134
rect 381062 621898 381146 622134
rect 381382 621898 381414 622134
rect 380794 582454 381414 621898
rect 380794 582218 380826 582454
rect 381062 582218 381146 582454
rect 381382 582218 381414 582454
rect 380794 582134 381414 582218
rect 380794 581898 380826 582134
rect 381062 581898 381146 582134
rect 381382 581898 381414 582134
rect 380794 542454 381414 581898
rect 380794 542218 380826 542454
rect 381062 542218 381146 542454
rect 381382 542218 381414 542454
rect 380794 542134 381414 542218
rect 380794 541898 380826 542134
rect 381062 541898 381146 542134
rect 381382 541898 381414 542134
rect 380794 502454 381414 541898
rect 380794 502218 380826 502454
rect 381062 502218 381146 502454
rect 381382 502218 381414 502454
rect 380794 502134 381414 502218
rect 380794 501898 380826 502134
rect 381062 501898 381146 502134
rect 381382 501898 381414 502134
rect 380794 462454 381414 501898
rect 380794 462218 380826 462454
rect 381062 462218 381146 462454
rect 381382 462218 381414 462454
rect 380794 462134 381414 462218
rect 380794 461898 380826 462134
rect 381062 461898 381146 462134
rect 381382 461898 381414 462134
rect 380794 422454 381414 461898
rect 380794 422218 380826 422454
rect 381062 422218 381146 422454
rect 381382 422218 381414 422454
rect 380794 422134 381414 422218
rect 380794 421898 380826 422134
rect 381062 421898 381146 422134
rect 381382 421898 381414 422134
rect 380794 382454 381414 421898
rect 380794 382218 380826 382454
rect 381062 382218 381146 382454
rect 381382 382218 381414 382454
rect 380794 382134 381414 382218
rect 380794 381898 380826 382134
rect 381062 381898 381146 382134
rect 381382 381898 381414 382134
rect 380794 342454 381414 381898
rect 380794 342218 380826 342454
rect 381062 342218 381146 342454
rect 381382 342218 381414 342454
rect 380794 342134 381414 342218
rect 380794 341898 380826 342134
rect 381062 341898 381146 342134
rect 381382 341898 381414 342134
rect 380794 302454 381414 341898
rect 380794 302218 380826 302454
rect 381062 302218 381146 302454
rect 381382 302218 381414 302454
rect 380794 302134 381414 302218
rect 380794 301898 380826 302134
rect 381062 301898 381146 302134
rect 381382 301898 381414 302134
rect 380794 262454 381414 301898
rect 380794 262218 380826 262454
rect 381062 262218 381146 262454
rect 381382 262218 381414 262454
rect 380794 262134 381414 262218
rect 380794 261898 380826 262134
rect 381062 261898 381146 262134
rect 381382 261898 381414 262134
rect 380794 222454 381414 261898
rect 380794 222218 380826 222454
rect 381062 222218 381146 222454
rect 381382 222218 381414 222454
rect 380794 222134 381414 222218
rect 380794 221898 380826 222134
rect 381062 221898 381146 222134
rect 381382 221898 381414 222134
rect 380794 182454 381414 221898
rect 380794 182218 380826 182454
rect 381062 182218 381146 182454
rect 381382 182218 381414 182454
rect 380794 182134 381414 182218
rect 380794 181898 380826 182134
rect 381062 181898 381146 182134
rect 381382 181898 381414 182134
rect 380794 142454 381414 181898
rect 380794 142218 380826 142454
rect 381062 142218 381146 142454
rect 381382 142218 381414 142454
rect 380794 142134 381414 142218
rect 380794 141898 380826 142134
rect 381062 141898 381146 142134
rect 381382 141898 381414 142134
rect 380794 102454 381414 141898
rect 380794 102218 380826 102454
rect 381062 102218 381146 102454
rect 381382 102218 381414 102454
rect 380794 102134 381414 102218
rect 380794 101898 380826 102134
rect 381062 101898 381146 102134
rect 381382 101898 381414 102134
rect 380794 62454 381414 101898
rect 380794 62218 380826 62454
rect 381062 62218 381146 62454
rect 381382 62218 381414 62454
rect 380794 62134 381414 62218
rect 380794 61898 380826 62134
rect 381062 61898 381146 62134
rect 381382 61898 381414 62134
rect 380794 22454 381414 61898
rect 380794 22218 380826 22454
rect 381062 22218 381146 22454
rect 381382 22218 381414 22454
rect 380794 22134 381414 22218
rect 380794 21898 380826 22134
rect 381062 21898 381146 22134
rect 381382 21898 381414 22134
rect 380794 -1306 381414 21898
rect 380794 -1542 380826 -1306
rect 381062 -1542 381146 -1306
rect 381382 -1542 381414 -1306
rect 380794 -1626 381414 -1542
rect 380794 -1862 380826 -1626
rect 381062 -1862 381146 -1626
rect 381382 -1862 381414 -1626
rect 380794 -1894 381414 -1862
rect 384514 666174 385134 707162
rect 384514 665938 384546 666174
rect 384782 665938 384866 666174
rect 385102 665938 385134 666174
rect 384514 665854 385134 665938
rect 384514 665618 384546 665854
rect 384782 665618 384866 665854
rect 385102 665618 385134 665854
rect 384514 626174 385134 665618
rect 384514 625938 384546 626174
rect 384782 625938 384866 626174
rect 385102 625938 385134 626174
rect 384514 625854 385134 625938
rect 384514 625618 384546 625854
rect 384782 625618 384866 625854
rect 385102 625618 385134 625854
rect 384514 586174 385134 625618
rect 384514 585938 384546 586174
rect 384782 585938 384866 586174
rect 385102 585938 385134 586174
rect 384514 585854 385134 585938
rect 384514 585618 384546 585854
rect 384782 585618 384866 585854
rect 385102 585618 385134 585854
rect 384514 546174 385134 585618
rect 384514 545938 384546 546174
rect 384782 545938 384866 546174
rect 385102 545938 385134 546174
rect 384514 545854 385134 545938
rect 384514 545618 384546 545854
rect 384782 545618 384866 545854
rect 385102 545618 385134 545854
rect 384514 506174 385134 545618
rect 384514 505938 384546 506174
rect 384782 505938 384866 506174
rect 385102 505938 385134 506174
rect 384514 505854 385134 505938
rect 384514 505618 384546 505854
rect 384782 505618 384866 505854
rect 385102 505618 385134 505854
rect 384514 466174 385134 505618
rect 384514 465938 384546 466174
rect 384782 465938 384866 466174
rect 385102 465938 385134 466174
rect 384514 465854 385134 465938
rect 384514 465618 384546 465854
rect 384782 465618 384866 465854
rect 385102 465618 385134 465854
rect 384514 426174 385134 465618
rect 384514 425938 384546 426174
rect 384782 425938 384866 426174
rect 385102 425938 385134 426174
rect 384514 425854 385134 425938
rect 384514 425618 384546 425854
rect 384782 425618 384866 425854
rect 385102 425618 385134 425854
rect 384514 386174 385134 425618
rect 384514 385938 384546 386174
rect 384782 385938 384866 386174
rect 385102 385938 385134 386174
rect 384514 385854 385134 385938
rect 384514 385618 384546 385854
rect 384782 385618 384866 385854
rect 385102 385618 385134 385854
rect 384514 346174 385134 385618
rect 384514 345938 384546 346174
rect 384782 345938 384866 346174
rect 385102 345938 385134 346174
rect 384514 345854 385134 345938
rect 384514 345618 384546 345854
rect 384782 345618 384866 345854
rect 385102 345618 385134 345854
rect 384514 306174 385134 345618
rect 384514 305938 384546 306174
rect 384782 305938 384866 306174
rect 385102 305938 385134 306174
rect 384514 305854 385134 305938
rect 384514 305618 384546 305854
rect 384782 305618 384866 305854
rect 385102 305618 385134 305854
rect 384514 266174 385134 305618
rect 384514 265938 384546 266174
rect 384782 265938 384866 266174
rect 385102 265938 385134 266174
rect 384514 265854 385134 265938
rect 384514 265618 384546 265854
rect 384782 265618 384866 265854
rect 385102 265618 385134 265854
rect 384514 226174 385134 265618
rect 384514 225938 384546 226174
rect 384782 225938 384866 226174
rect 385102 225938 385134 226174
rect 384514 225854 385134 225938
rect 384514 225618 384546 225854
rect 384782 225618 384866 225854
rect 385102 225618 385134 225854
rect 384514 186174 385134 225618
rect 384514 185938 384546 186174
rect 384782 185938 384866 186174
rect 385102 185938 385134 186174
rect 384514 185854 385134 185938
rect 384514 185618 384546 185854
rect 384782 185618 384866 185854
rect 385102 185618 385134 185854
rect 384514 146174 385134 185618
rect 384514 145938 384546 146174
rect 384782 145938 384866 146174
rect 385102 145938 385134 146174
rect 384514 145854 385134 145938
rect 384514 145618 384546 145854
rect 384782 145618 384866 145854
rect 385102 145618 385134 145854
rect 384514 106174 385134 145618
rect 384514 105938 384546 106174
rect 384782 105938 384866 106174
rect 385102 105938 385134 106174
rect 384514 105854 385134 105938
rect 384514 105618 384546 105854
rect 384782 105618 384866 105854
rect 385102 105618 385134 105854
rect 384514 66174 385134 105618
rect 384514 65938 384546 66174
rect 384782 65938 384866 66174
rect 385102 65938 385134 66174
rect 384514 65854 385134 65938
rect 384514 65618 384546 65854
rect 384782 65618 384866 65854
rect 385102 65618 385134 65854
rect 384514 26174 385134 65618
rect 384514 25938 384546 26174
rect 384782 25938 384866 26174
rect 385102 25938 385134 26174
rect 384514 25854 385134 25938
rect 384514 25618 384546 25854
rect 384782 25618 384866 25854
rect 385102 25618 385134 25854
rect 384514 -3226 385134 25618
rect 384514 -3462 384546 -3226
rect 384782 -3462 384866 -3226
rect 385102 -3462 385134 -3226
rect 384514 -3546 385134 -3462
rect 384514 -3782 384546 -3546
rect 384782 -3782 384866 -3546
rect 385102 -3782 385134 -3546
rect 384514 -3814 385134 -3782
rect 388234 669894 388854 709082
rect 388234 669658 388266 669894
rect 388502 669658 388586 669894
rect 388822 669658 388854 669894
rect 388234 669574 388854 669658
rect 388234 669338 388266 669574
rect 388502 669338 388586 669574
rect 388822 669338 388854 669574
rect 388234 629894 388854 669338
rect 388234 629658 388266 629894
rect 388502 629658 388586 629894
rect 388822 629658 388854 629894
rect 388234 629574 388854 629658
rect 388234 629338 388266 629574
rect 388502 629338 388586 629574
rect 388822 629338 388854 629574
rect 388234 589894 388854 629338
rect 388234 589658 388266 589894
rect 388502 589658 388586 589894
rect 388822 589658 388854 589894
rect 388234 589574 388854 589658
rect 388234 589338 388266 589574
rect 388502 589338 388586 589574
rect 388822 589338 388854 589574
rect 388234 549894 388854 589338
rect 388234 549658 388266 549894
rect 388502 549658 388586 549894
rect 388822 549658 388854 549894
rect 388234 549574 388854 549658
rect 388234 549338 388266 549574
rect 388502 549338 388586 549574
rect 388822 549338 388854 549574
rect 388234 509894 388854 549338
rect 388234 509658 388266 509894
rect 388502 509658 388586 509894
rect 388822 509658 388854 509894
rect 388234 509574 388854 509658
rect 388234 509338 388266 509574
rect 388502 509338 388586 509574
rect 388822 509338 388854 509574
rect 388234 469894 388854 509338
rect 388234 469658 388266 469894
rect 388502 469658 388586 469894
rect 388822 469658 388854 469894
rect 388234 469574 388854 469658
rect 388234 469338 388266 469574
rect 388502 469338 388586 469574
rect 388822 469338 388854 469574
rect 388234 429894 388854 469338
rect 388234 429658 388266 429894
rect 388502 429658 388586 429894
rect 388822 429658 388854 429894
rect 388234 429574 388854 429658
rect 388234 429338 388266 429574
rect 388502 429338 388586 429574
rect 388822 429338 388854 429574
rect 388234 389894 388854 429338
rect 388234 389658 388266 389894
rect 388502 389658 388586 389894
rect 388822 389658 388854 389894
rect 388234 389574 388854 389658
rect 388234 389338 388266 389574
rect 388502 389338 388586 389574
rect 388822 389338 388854 389574
rect 388234 349894 388854 389338
rect 388234 349658 388266 349894
rect 388502 349658 388586 349894
rect 388822 349658 388854 349894
rect 388234 349574 388854 349658
rect 388234 349338 388266 349574
rect 388502 349338 388586 349574
rect 388822 349338 388854 349574
rect 388234 309894 388854 349338
rect 388234 309658 388266 309894
rect 388502 309658 388586 309894
rect 388822 309658 388854 309894
rect 388234 309574 388854 309658
rect 388234 309338 388266 309574
rect 388502 309338 388586 309574
rect 388822 309338 388854 309574
rect 388234 269894 388854 309338
rect 388234 269658 388266 269894
rect 388502 269658 388586 269894
rect 388822 269658 388854 269894
rect 388234 269574 388854 269658
rect 388234 269338 388266 269574
rect 388502 269338 388586 269574
rect 388822 269338 388854 269574
rect 388234 229894 388854 269338
rect 388234 229658 388266 229894
rect 388502 229658 388586 229894
rect 388822 229658 388854 229894
rect 388234 229574 388854 229658
rect 388234 229338 388266 229574
rect 388502 229338 388586 229574
rect 388822 229338 388854 229574
rect 388234 189894 388854 229338
rect 388234 189658 388266 189894
rect 388502 189658 388586 189894
rect 388822 189658 388854 189894
rect 388234 189574 388854 189658
rect 388234 189338 388266 189574
rect 388502 189338 388586 189574
rect 388822 189338 388854 189574
rect 388234 149894 388854 189338
rect 388234 149658 388266 149894
rect 388502 149658 388586 149894
rect 388822 149658 388854 149894
rect 388234 149574 388854 149658
rect 388234 149338 388266 149574
rect 388502 149338 388586 149574
rect 388822 149338 388854 149574
rect 388234 109894 388854 149338
rect 388234 109658 388266 109894
rect 388502 109658 388586 109894
rect 388822 109658 388854 109894
rect 388234 109574 388854 109658
rect 388234 109338 388266 109574
rect 388502 109338 388586 109574
rect 388822 109338 388854 109574
rect 388234 69894 388854 109338
rect 388234 69658 388266 69894
rect 388502 69658 388586 69894
rect 388822 69658 388854 69894
rect 388234 69574 388854 69658
rect 388234 69338 388266 69574
rect 388502 69338 388586 69574
rect 388822 69338 388854 69574
rect 388234 29894 388854 69338
rect 388234 29658 388266 29894
rect 388502 29658 388586 29894
rect 388822 29658 388854 29894
rect 388234 29574 388854 29658
rect 388234 29338 388266 29574
rect 388502 29338 388586 29574
rect 388822 29338 388854 29574
rect 388234 -5146 388854 29338
rect 388234 -5382 388266 -5146
rect 388502 -5382 388586 -5146
rect 388822 -5382 388854 -5146
rect 388234 -5466 388854 -5382
rect 388234 -5702 388266 -5466
rect 388502 -5702 388586 -5466
rect 388822 -5702 388854 -5466
rect 388234 -5734 388854 -5702
rect 391954 673614 392574 711002
rect 411954 710598 412574 711590
rect 411954 710362 411986 710598
rect 412222 710362 412306 710598
rect 412542 710362 412574 710598
rect 411954 710278 412574 710362
rect 411954 710042 411986 710278
rect 412222 710042 412306 710278
rect 412542 710042 412574 710278
rect 408234 708678 408854 709670
rect 408234 708442 408266 708678
rect 408502 708442 408586 708678
rect 408822 708442 408854 708678
rect 408234 708358 408854 708442
rect 408234 708122 408266 708358
rect 408502 708122 408586 708358
rect 408822 708122 408854 708358
rect 404514 706758 405134 707750
rect 404514 706522 404546 706758
rect 404782 706522 404866 706758
rect 405102 706522 405134 706758
rect 404514 706438 405134 706522
rect 404514 706202 404546 706438
rect 404782 706202 404866 706438
rect 405102 706202 405134 706438
rect 391954 673378 391986 673614
rect 392222 673378 392306 673614
rect 392542 673378 392574 673614
rect 391954 673294 392574 673378
rect 391954 673058 391986 673294
rect 392222 673058 392306 673294
rect 392542 673058 392574 673294
rect 391954 633614 392574 673058
rect 391954 633378 391986 633614
rect 392222 633378 392306 633614
rect 392542 633378 392574 633614
rect 391954 633294 392574 633378
rect 391954 633058 391986 633294
rect 392222 633058 392306 633294
rect 392542 633058 392574 633294
rect 391954 593614 392574 633058
rect 391954 593378 391986 593614
rect 392222 593378 392306 593614
rect 392542 593378 392574 593614
rect 391954 593294 392574 593378
rect 391954 593058 391986 593294
rect 392222 593058 392306 593294
rect 392542 593058 392574 593294
rect 391954 553614 392574 593058
rect 391954 553378 391986 553614
rect 392222 553378 392306 553614
rect 392542 553378 392574 553614
rect 391954 553294 392574 553378
rect 391954 553058 391986 553294
rect 392222 553058 392306 553294
rect 392542 553058 392574 553294
rect 391954 513614 392574 553058
rect 391954 513378 391986 513614
rect 392222 513378 392306 513614
rect 392542 513378 392574 513614
rect 391954 513294 392574 513378
rect 391954 513058 391986 513294
rect 392222 513058 392306 513294
rect 392542 513058 392574 513294
rect 391954 473614 392574 513058
rect 391954 473378 391986 473614
rect 392222 473378 392306 473614
rect 392542 473378 392574 473614
rect 391954 473294 392574 473378
rect 391954 473058 391986 473294
rect 392222 473058 392306 473294
rect 392542 473058 392574 473294
rect 391954 433614 392574 473058
rect 391954 433378 391986 433614
rect 392222 433378 392306 433614
rect 392542 433378 392574 433614
rect 391954 433294 392574 433378
rect 391954 433058 391986 433294
rect 392222 433058 392306 433294
rect 392542 433058 392574 433294
rect 391954 393614 392574 433058
rect 391954 393378 391986 393614
rect 392222 393378 392306 393614
rect 392542 393378 392574 393614
rect 391954 393294 392574 393378
rect 391954 393058 391986 393294
rect 392222 393058 392306 393294
rect 392542 393058 392574 393294
rect 391954 353614 392574 393058
rect 391954 353378 391986 353614
rect 392222 353378 392306 353614
rect 392542 353378 392574 353614
rect 391954 353294 392574 353378
rect 391954 353058 391986 353294
rect 392222 353058 392306 353294
rect 392542 353058 392574 353294
rect 391954 313614 392574 353058
rect 391954 313378 391986 313614
rect 392222 313378 392306 313614
rect 392542 313378 392574 313614
rect 391954 313294 392574 313378
rect 391954 313058 391986 313294
rect 392222 313058 392306 313294
rect 392542 313058 392574 313294
rect 391954 273614 392574 313058
rect 391954 273378 391986 273614
rect 392222 273378 392306 273614
rect 392542 273378 392574 273614
rect 391954 273294 392574 273378
rect 391954 273058 391986 273294
rect 392222 273058 392306 273294
rect 392542 273058 392574 273294
rect 391954 233614 392574 273058
rect 391954 233378 391986 233614
rect 392222 233378 392306 233614
rect 392542 233378 392574 233614
rect 391954 233294 392574 233378
rect 391954 233058 391986 233294
rect 392222 233058 392306 233294
rect 392542 233058 392574 233294
rect 391954 193614 392574 233058
rect 391954 193378 391986 193614
rect 392222 193378 392306 193614
rect 392542 193378 392574 193614
rect 391954 193294 392574 193378
rect 391954 193058 391986 193294
rect 392222 193058 392306 193294
rect 392542 193058 392574 193294
rect 391954 153614 392574 193058
rect 391954 153378 391986 153614
rect 392222 153378 392306 153614
rect 392542 153378 392574 153614
rect 391954 153294 392574 153378
rect 391954 153058 391986 153294
rect 392222 153058 392306 153294
rect 392542 153058 392574 153294
rect 391954 113614 392574 153058
rect 391954 113378 391986 113614
rect 392222 113378 392306 113614
rect 392542 113378 392574 113614
rect 391954 113294 392574 113378
rect 391954 113058 391986 113294
rect 392222 113058 392306 113294
rect 392542 113058 392574 113294
rect 391954 73614 392574 113058
rect 391954 73378 391986 73614
rect 392222 73378 392306 73614
rect 392542 73378 392574 73614
rect 391954 73294 392574 73378
rect 391954 73058 391986 73294
rect 392222 73058 392306 73294
rect 392542 73058 392574 73294
rect 391954 33614 392574 73058
rect 391954 33378 391986 33614
rect 392222 33378 392306 33614
rect 392542 33378 392574 33614
rect 391954 33294 392574 33378
rect 391954 33058 391986 33294
rect 392222 33058 392306 33294
rect 392542 33058 392574 33294
rect 371954 -6342 371986 -6106
rect 372222 -6342 372306 -6106
rect 372542 -6342 372574 -6106
rect 371954 -6426 372574 -6342
rect 371954 -6662 371986 -6426
rect 372222 -6662 372306 -6426
rect 372542 -6662 372574 -6426
rect 371954 -7654 372574 -6662
rect 391954 -7066 392574 33058
rect 400794 704838 401414 705830
rect 400794 704602 400826 704838
rect 401062 704602 401146 704838
rect 401382 704602 401414 704838
rect 400794 704518 401414 704602
rect 400794 704282 400826 704518
rect 401062 704282 401146 704518
rect 401382 704282 401414 704518
rect 400794 682454 401414 704282
rect 400794 682218 400826 682454
rect 401062 682218 401146 682454
rect 401382 682218 401414 682454
rect 400794 682134 401414 682218
rect 400794 681898 400826 682134
rect 401062 681898 401146 682134
rect 401382 681898 401414 682134
rect 400794 642454 401414 681898
rect 400794 642218 400826 642454
rect 401062 642218 401146 642454
rect 401382 642218 401414 642454
rect 400794 642134 401414 642218
rect 400794 641898 400826 642134
rect 401062 641898 401146 642134
rect 401382 641898 401414 642134
rect 400794 602454 401414 641898
rect 400794 602218 400826 602454
rect 401062 602218 401146 602454
rect 401382 602218 401414 602454
rect 400794 602134 401414 602218
rect 400794 601898 400826 602134
rect 401062 601898 401146 602134
rect 401382 601898 401414 602134
rect 400794 562454 401414 601898
rect 400794 562218 400826 562454
rect 401062 562218 401146 562454
rect 401382 562218 401414 562454
rect 400794 562134 401414 562218
rect 400794 561898 400826 562134
rect 401062 561898 401146 562134
rect 401382 561898 401414 562134
rect 400794 522454 401414 561898
rect 400794 522218 400826 522454
rect 401062 522218 401146 522454
rect 401382 522218 401414 522454
rect 400794 522134 401414 522218
rect 400794 521898 400826 522134
rect 401062 521898 401146 522134
rect 401382 521898 401414 522134
rect 400794 482454 401414 521898
rect 400794 482218 400826 482454
rect 401062 482218 401146 482454
rect 401382 482218 401414 482454
rect 400794 482134 401414 482218
rect 400794 481898 400826 482134
rect 401062 481898 401146 482134
rect 401382 481898 401414 482134
rect 400794 442454 401414 481898
rect 400794 442218 400826 442454
rect 401062 442218 401146 442454
rect 401382 442218 401414 442454
rect 400794 442134 401414 442218
rect 400794 441898 400826 442134
rect 401062 441898 401146 442134
rect 401382 441898 401414 442134
rect 400794 402454 401414 441898
rect 400794 402218 400826 402454
rect 401062 402218 401146 402454
rect 401382 402218 401414 402454
rect 400794 402134 401414 402218
rect 400794 401898 400826 402134
rect 401062 401898 401146 402134
rect 401382 401898 401414 402134
rect 400794 362454 401414 401898
rect 400794 362218 400826 362454
rect 401062 362218 401146 362454
rect 401382 362218 401414 362454
rect 400794 362134 401414 362218
rect 400794 361898 400826 362134
rect 401062 361898 401146 362134
rect 401382 361898 401414 362134
rect 400794 322454 401414 361898
rect 400794 322218 400826 322454
rect 401062 322218 401146 322454
rect 401382 322218 401414 322454
rect 400794 322134 401414 322218
rect 400794 321898 400826 322134
rect 401062 321898 401146 322134
rect 401382 321898 401414 322134
rect 400794 282454 401414 321898
rect 400794 282218 400826 282454
rect 401062 282218 401146 282454
rect 401382 282218 401414 282454
rect 400794 282134 401414 282218
rect 400794 281898 400826 282134
rect 401062 281898 401146 282134
rect 401382 281898 401414 282134
rect 400794 242454 401414 281898
rect 400794 242218 400826 242454
rect 401062 242218 401146 242454
rect 401382 242218 401414 242454
rect 400794 242134 401414 242218
rect 400794 241898 400826 242134
rect 401062 241898 401146 242134
rect 401382 241898 401414 242134
rect 400794 202454 401414 241898
rect 400794 202218 400826 202454
rect 401062 202218 401146 202454
rect 401382 202218 401414 202454
rect 400794 202134 401414 202218
rect 400794 201898 400826 202134
rect 401062 201898 401146 202134
rect 401382 201898 401414 202134
rect 400794 162454 401414 201898
rect 400794 162218 400826 162454
rect 401062 162218 401146 162454
rect 401382 162218 401414 162454
rect 400794 162134 401414 162218
rect 400794 161898 400826 162134
rect 401062 161898 401146 162134
rect 401382 161898 401414 162134
rect 400794 122454 401414 161898
rect 400794 122218 400826 122454
rect 401062 122218 401146 122454
rect 401382 122218 401414 122454
rect 400794 122134 401414 122218
rect 400794 121898 400826 122134
rect 401062 121898 401146 122134
rect 401382 121898 401414 122134
rect 400794 82454 401414 121898
rect 400794 82218 400826 82454
rect 401062 82218 401146 82454
rect 401382 82218 401414 82454
rect 400794 82134 401414 82218
rect 400794 81898 400826 82134
rect 401062 81898 401146 82134
rect 401382 81898 401414 82134
rect 400794 42454 401414 81898
rect 400794 42218 400826 42454
rect 401062 42218 401146 42454
rect 401382 42218 401414 42454
rect 400794 42134 401414 42218
rect 400794 41898 400826 42134
rect 401062 41898 401146 42134
rect 401382 41898 401414 42134
rect 400794 2454 401414 41898
rect 400794 2218 400826 2454
rect 401062 2218 401146 2454
rect 401382 2218 401414 2454
rect 400794 2134 401414 2218
rect 400794 1898 400826 2134
rect 401062 1898 401146 2134
rect 401382 1898 401414 2134
rect 400794 -346 401414 1898
rect 400794 -582 400826 -346
rect 401062 -582 401146 -346
rect 401382 -582 401414 -346
rect 400794 -666 401414 -582
rect 400794 -902 400826 -666
rect 401062 -902 401146 -666
rect 401382 -902 401414 -666
rect 400794 -1894 401414 -902
rect 404514 686174 405134 706202
rect 404514 685938 404546 686174
rect 404782 685938 404866 686174
rect 405102 685938 405134 686174
rect 404514 685854 405134 685938
rect 404514 685618 404546 685854
rect 404782 685618 404866 685854
rect 405102 685618 405134 685854
rect 404514 646174 405134 685618
rect 404514 645938 404546 646174
rect 404782 645938 404866 646174
rect 405102 645938 405134 646174
rect 404514 645854 405134 645938
rect 404514 645618 404546 645854
rect 404782 645618 404866 645854
rect 405102 645618 405134 645854
rect 404514 606174 405134 645618
rect 404514 605938 404546 606174
rect 404782 605938 404866 606174
rect 405102 605938 405134 606174
rect 404514 605854 405134 605938
rect 404514 605618 404546 605854
rect 404782 605618 404866 605854
rect 405102 605618 405134 605854
rect 404514 566174 405134 605618
rect 404514 565938 404546 566174
rect 404782 565938 404866 566174
rect 405102 565938 405134 566174
rect 404514 565854 405134 565938
rect 404514 565618 404546 565854
rect 404782 565618 404866 565854
rect 405102 565618 405134 565854
rect 404514 526174 405134 565618
rect 404514 525938 404546 526174
rect 404782 525938 404866 526174
rect 405102 525938 405134 526174
rect 404514 525854 405134 525938
rect 404514 525618 404546 525854
rect 404782 525618 404866 525854
rect 405102 525618 405134 525854
rect 404514 486174 405134 525618
rect 404514 485938 404546 486174
rect 404782 485938 404866 486174
rect 405102 485938 405134 486174
rect 404514 485854 405134 485938
rect 404514 485618 404546 485854
rect 404782 485618 404866 485854
rect 405102 485618 405134 485854
rect 404514 446174 405134 485618
rect 404514 445938 404546 446174
rect 404782 445938 404866 446174
rect 405102 445938 405134 446174
rect 404514 445854 405134 445938
rect 404514 445618 404546 445854
rect 404782 445618 404866 445854
rect 405102 445618 405134 445854
rect 404514 406174 405134 445618
rect 404514 405938 404546 406174
rect 404782 405938 404866 406174
rect 405102 405938 405134 406174
rect 404514 405854 405134 405938
rect 404514 405618 404546 405854
rect 404782 405618 404866 405854
rect 405102 405618 405134 405854
rect 404514 366174 405134 405618
rect 404514 365938 404546 366174
rect 404782 365938 404866 366174
rect 405102 365938 405134 366174
rect 404514 365854 405134 365938
rect 404514 365618 404546 365854
rect 404782 365618 404866 365854
rect 405102 365618 405134 365854
rect 404514 326174 405134 365618
rect 404514 325938 404546 326174
rect 404782 325938 404866 326174
rect 405102 325938 405134 326174
rect 404514 325854 405134 325938
rect 404514 325618 404546 325854
rect 404782 325618 404866 325854
rect 405102 325618 405134 325854
rect 404514 286174 405134 325618
rect 404514 285938 404546 286174
rect 404782 285938 404866 286174
rect 405102 285938 405134 286174
rect 404514 285854 405134 285938
rect 404514 285618 404546 285854
rect 404782 285618 404866 285854
rect 405102 285618 405134 285854
rect 404514 246174 405134 285618
rect 404514 245938 404546 246174
rect 404782 245938 404866 246174
rect 405102 245938 405134 246174
rect 404514 245854 405134 245938
rect 404514 245618 404546 245854
rect 404782 245618 404866 245854
rect 405102 245618 405134 245854
rect 404514 206174 405134 245618
rect 404514 205938 404546 206174
rect 404782 205938 404866 206174
rect 405102 205938 405134 206174
rect 404514 205854 405134 205938
rect 404514 205618 404546 205854
rect 404782 205618 404866 205854
rect 405102 205618 405134 205854
rect 404514 166174 405134 205618
rect 404514 165938 404546 166174
rect 404782 165938 404866 166174
rect 405102 165938 405134 166174
rect 404514 165854 405134 165938
rect 404514 165618 404546 165854
rect 404782 165618 404866 165854
rect 405102 165618 405134 165854
rect 404514 126174 405134 165618
rect 404514 125938 404546 126174
rect 404782 125938 404866 126174
rect 405102 125938 405134 126174
rect 404514 125854 405134 125938
rect 404514 125618 404546 125854
rect 404782 125618 404866 125854
rect 405102 125618 405134 125854
rect 404514 86174 405134 125618
rect 404514 85938 404546 86174
rect 404782 85938 404866 86174
rect 405102 85938 405134 86174
rect 404514 85854 405134 85938
rect 404514 85618 404546 85854
rect 404782 85618 404866 85854
rect 405102 85618 405134 85854
rect 404514 46174 405134 85618
rect 404514 45938 404546 46174
rect 404782 45938 404866 46174
rect 405102 45938 405134 46174
rect 404514 45854 405134 45938
rect 404514 45618 404546 45854
rect 404782 45618 404866 45854
rect 405102 45618 405134 45854
rect 404514 6174 405134 45618
rect 404514 5938 404546 6174
rect 404782 5938 404866 6174
rect 405102 5938 405134 6174
rect 404514 5854 405134 5938
rect 404514 5618 404546 5854
rect 404782 5618 404866 5854
rect 405102 5618 405134 5854
rect 404514 -2266 405134 5618
rect 404514 -2502 404546 -2266
rect 404782 -2502 404866 -2266
rect 405102 -2502 405134 -2266
rect 404514 -2586 405134 -2502
rect 404514 -2822 404546 -2586
rect 404782 -2822 404866 -2586
rect 405102 -2822 405134 -2586
rect 404514 -3814 405134 -2822
rect 408234 689894 408854 708122
rect 408234 689658 408266 689894
rect 408502 689658 408586 689894
rect 408822 689658 408854 689894
rect 408234 689574 408854 689658
rect 408234 689338 408266 689574
rect 408502 689338 408586 689574
rect 408822 689338 408854 689574
rect 408234 649894 408854 689338
rect 408234 649658 408266 649894
rect 408502 649658 408586 649894
rect 408822 649658 408854 649894
rect 408234 649574 408854 649658
rect 408234 649338 408266 649574
rect 408502 649338 408586 649574
rect 408822 649338 408854 649574
rect 408234 609894 408854 649338
rect 408234 609658 408266 609894
rect 408502 609658 408586 609894
rect 408822 609658 408854 609894
rect 408234 609574 408854 609658
rect 408234 609338 408266 609574
rect 408502 609338 408586 609574
rect 408822 609338 408854 609574
rect 408234 569894 408854 609338
rect 408234 569658 408266 569894
rect 408502 569658 408586 569894
rect 408822 569658 408854 569894
rect 408234 569574 408854 569658
rect 408234 569338 408266 569574
rect 408502 569338 408586 569574
rect 408822 569338 408854 569574
rect 408234 529894 408854 569338
rect 408234 529658 408266 529894
rect 408502 529658 408586 529894
rect 408822 529658 408854 529894
rect 408234 529574 408854 529658
rect 408234 529338 408266 529574
rect 408502 529338 408586 529574
rect 408822 529338 408854 529574
rect 408234 489894 408854 529338
rect 408234 489658 408266 489894
rect 408502 489658 408586 489894
rect 408822 489658 408854 489894
rect 408234 489574 408854 489658
rect 408234 489338 408266 489574
rect 408502 489338 408586 489574
rect 408822 489338 408854 489574
rect 408234 449894 408854 489338
rect 408234 449658 408266 449894
rect 408502 449658 408586 449894
rect 408822 449658 408854 449894
rect 408234 449574 408854 449658
rect 408234 449338 408266 449574
rect 408502 449338 408586 449574
rect 408822 449338 408854 449574
rect 408234 409894 408854 449338
rect 408234 409658 408266 409894
rect 408502 409658 408586 409894
rect 408822 409658 408854 409894
rect 408234 409574 408854 409658
rect 408234 409338 408266 409574
rect 408502 409338 408586 409574
rect 408822 409338 408854 409574
rect 408234 369894 408854 409338
rect 408234 369658 408266 369894
rect 408502 369658 408586 369894
rect 408822 369658 408854 369894
rect 408234 369574 408854 369658
rect 408234 369338 408266 369574
rect 408502 369338 408586 369574
rect 408822 369338 408854 369574
rect 408234 329894 408854 369338
rect 408234 329658 408266 329894
rect 408502 329658 408586 329894
rect 408822 329658 408854 329894
rect 408234 329574 408854 329658
rect 408234 329338 408266 329574
rect 408502 329338 408586 329574
rect 408822 329338 408854 329574
rect 408234 289894 408854 329338
rect 408234 289658 408266 289894
rect 408502 289658 408586 289894
rect 408822 289658 408854 289894
rect 408234 289574 408854 289658
rect 408234 289338 408266 289574
rect 408502 289338 408586 289574
rect 408822 289338 408854 289574
rect 408234 249894 408854 289338
rect 408234 249658 408266 249894
rect 408502 249658 408586 249894
rect 408822 249658 408854 249894
rect 408234 249574 408854 249658
rect 408234 249338 408266 249574
rect 408502 249338 408586 249574
rect 408822 249338 408854 249574
rect 408234 209894 408854 249338
rect 408234 209658 408266 209894
rect 408502 209658 408586 209894
rect 408822 209658 408854 209894
rect 408234 209574 408854 209658
rect 408234 209338 408266 209574
rect 408502 209338 408586 209574
rect 408822 209338 408854 209574
rect 408234 169894 408854 209338
rect 408234 169658 408266 169894
rect 408502 169658 408586 169894
rect 408822 169658 408854 169894
rect 408234 169574 408854 169658
rect 408234 169338 408266 169574
rect 408502 169338 408586 169574
rect 408822 169338 408854 169574
rect 408234 129894 408854 169338
rect 408234 129658 408266 129894
rect 408502 129658 408586 129894
rect 408822 129658 408854 129894
rect 408234 129574 408854 129658
rect 408234 129338 408266 129574
rect 408502 129338 408586 129574
rect 408822 129338 408854 129574
rect 408234 89894 408854 129338
rect 408234 89658 408266 89894
rect 408502 89658 408586 89894
rect 408822 89658 408854 89894
rect 408234 89574 408854 89658
rect 408234 89338 408266 89574
rect 408502 89338 408586 89574
rect 408822 89338 408854 89574
rect 408234 49894 408854 89338
rect 408234 49658 408266 49894
rect 408502 49658 408586 49894
rect 408822 49658 408854 49894
rect 408234 49574 408854 49658
rect 408234 49338 408266 49574
rect 408502 49338 408586 49574
rect 408822 49338 408854 49574
rect 408234 9894 408854 49338
rect 408234 9658 408266 9894
rect 408502 9658 408586 9894
rect 408822 9658 408854 9894
rect 408234 9574 408854 9658
rect 408234 9338 408266 9574
rect 408502 9338 408586 9574
rect 408822 9338 408854 9574
rect 408234 -4186 408854 9338
rect 408234 -4422 408266 -4186
rect 408502 -4422 408586 -4186
rect 408822 -4422 408854 -4186
rect 408234 -4506 408854 -4422
rect 408234 -4742 408266 -4506
rect 408502 -4742 408586 -4506
rect 408822 -4742 408854 -4506
rect 408234 -5734 408854 -4742
rect 411954 693614 412574 710042
rect 431954 711558 432574 711590
rect 431954 711322 431986 711558
rect 432222 711322 432306 711558
rect 432542 711322 432574 711558
rect 431954 711238 432574 711322
rect 431954 711002 431986 711238
rect 432222 711002 432306 711238
rect 432542 711002 432574 711238
rect 428234 709638 428854 709670
rect 428234 709402 428266 709638
rect 428502 709402 428586 709638
rect 428822 709402 428854 709638
rect 428234 709318 428854 709402
rect 428234 709082 428266 709318
rect 428502 709082 428586 709318
rect 428822 709082 428854 709318
rect 424514 707718 425134 707750
rect 424514 707482 424546 707718
rect 424782 707482 424866 707718
rect 425102 707482 425134 707718
rect 424514 707398 425134 707482
rect 424514 707162 424546 707398
rect 424782 707162 424866 707398
rect 425102 707162 425134 707398
rect 411954 693378 411986 693614
rect 412222 693378 412306 693614
rect 412542 693378 412574 693614
rect 411954 693294 412574 693378
rect 411954 693058 411986 693294
rect 412222 693058 412306 693294
rect 412542 693058 412574 693294
rect 411954 653614 412574 693058
rect 411954 653378 411986 653614
rect 412222 653378 412306 653614
rect 412542 653378 412574 653614
rect 411954 653294 412574 653378
rect 411954 653058 411986 653294
rect 412222 653058 412306 653294
rect 412542 653058 412574 653294
rect 411954 613614 412574 653058
rect 411954 613378 411986 613614
rect 412222 613378 412306 613614
rect 412542 613378 412574 613614
rect 411954 613294 412574 613378
rect 411954 613058 411986 613294
rect 412222 613058 412306 613294
rect 412542 613058 412574 613294
rect 411954 573614 412574 613058
rect 411954 573378 411986 573614
rect 412222 573378 412306 573614
rect 412542 573378 412574 573614
rect 411954 573294 412574 573378
rect 411954 573058 411986 573294
rect 412222 573058 412306 573294
rect 412542 573058 412574 573294
rect 411954 533614 412574 573058
rect 411954 533378 411986 533614
rect 412222 533378 412306 533614
rect 412542 533378 412574 533614
rect 411954 533294 412574 533378
rect 411954 533058 411986 533294
rect 412222 533058 412306 533294
rect 412542 533058 412574 533294
rect 411954 493614 412574 533058
rect 411954 493378 411986 493614
rect 412222 493378 412306 493614
rect 412542 493378 412574 493614
rect 411954 493294 412574 493378
rect 411954 493058 411986 493294
rect 412222 493058 412306 493294
rect 412542 493058 412574 493294
rect 411954 453614 412574 493058
rect 411954 453378 411986 453614
rect 412222 453378 412306 453614
rect 412542 453378 412574 453614
rect 411954 453294 412574 453378
rect 411954 453058 411986 453294
rect 412222 453058 412306 453294
rect 412542 453058 412574 453294
rect 411954 413614 412574 453058
rect 411954 413378 411986 413614
rect 412222 413378 412306 413614
rect 412542 413378 412574 413614
rect 411954 413294 412574 413378
rect 411954 413058 411986 413294
rect 412222 413058 412306 413294
rect 412542 413058 412574 413294
rect 411954 373614 412574 413058
rect 411954 373378 411986 373614
rect 412222 373378 412306 373614
rect 412542 373378 412574 373614
rect 411954 373294 412574 373378
rect 411954 373058 411986 373294
rect 412222 373058 412306 373294
rect 412542 373058 412574 373294
rect 411954 333614 412574 373058
rect 411954 333378 411986 333614
rect 412222 333378 412306 333614
rect 412542 333378 412574 333614
rect 411954 333294 412574 333378
rect 411954 333058 411986 333294
rect 412222 333058 412306 333294
rect 412542 333058 412574 333294
rect 411954 293614 412574 333058
rect 411954 293378 411986 293614
rect 412222 293378 412306 293614
rect 412542 293378 412574 293614
rect 411954 293294 412574 293378
rect 411954 293058 411986 293294
rect 412222 293058 412306 293294
rect 412542 293058 412574 293294
rect 411954 253614 412574 293058
rect 411954 253378 411986 253614
rect 412222 253378 412306 253614
rect 412542 253378 412574 253614
rect 411954 253294 412574 253378
rect 411954 253058 411986 253294
rect 412222 253058 412306 253294
rect 412542 253058 412574 253294
rect 411954 213614 412574 253058
rect 411954 213378 411986 213614
rect 412222 213378 412306 213614
rect 412542 213378 412574 213614
rect 411954 213294 412574 213378
rect 411954 213058 411986 213294
rect 412222 213058 412306 213294
rect 412542 213058 412574 213294
rect 411954 173614 412574 213058
rect 411954 173378 411986 173614
rect 412222 173378 412306 173614
rect 412542 173378 412574 173614
rect 411954 173294 412574 173378
rect 411954 173058 411986 173294
rect 412222 173058 412306 173294
rect 412542 173058 412574 173294
rect 411954 133614 412574 173058
rect 411954 133378 411986 133614
rect 412222 133378 412306 133614
rect 412542 133378 412574 133614
rect 411954 133294 412574 133378
rect 411954 133058 411986 133294
rect 412222 133058 412306 133294
rect 412542 133058 412574 133294
rect 411954 93614 412574 133058
rect 411954 93378 411986 93614
rect 412222 93378 412306 93614
rect 412542 93378 412574 93614
rect 411954 93294 412574 93378
rect 411954 93058 411986 93294
rect 412222 93058 412306 93294
rect 412542 93058 412574 93294
rect 411954 53614 412574 93058
rect 411954 53378 411986 53614
rect 412222 53378 412306 53614
rect 412542 53378 412574 53614
rect 411954 53294 412574 53378
rect 411954 53058 411986 53294
rect 412222 53058 412306 53294
rect 412542 53058 412574 53294
rect 411954 13614 412574 53058
rect 411954 13378 411986 13614
rect 412222 13378 412306 13614
rect 412542 13378 412574 13614
rect 411954 13294 412574 13378
rect 411954 13058 411986 13294
rect 412222 13058 412306 13294
rect 412542 13058 412574 13294
rect 391954 -7302 391986 -7066
rect 392222 -7302 392306 -7066
rect 392542 -7302 392574 -7066
rect 391954 -7386 392574 -7302
rect 391954 -7622 391986 -7386
rect 392222 -7622 392306 -7386
rect 392542 -7622 392574 -7386
rect 391954 -7654 392574 -7622
rect 411954 -6106 412574 13058
rect 420794 705798 421414 705830
rect 420794 705562 420826 705798
rect 421062 705562 421146 705798
rect 421382 705562 421414 705798
rect 420794 705478 421414 705562
rect 420794 705242 420826 705478
rect 421062 705242 421146 705478
rect 421382 705242 421414 705478
rect 420794 662454 421414 705242
rect 420794 662218 420826 662454
rect 421062 662218 421146 662454
rect 421382 662218 421414 662454
rect 420794 662134 421414 662218
rect 420794 661898 420826 662134
rect 421062 661898 421146 662134
rect 421382 661898 421414 662134
rect 420794 622454 421414 661898
rect 420794 622218 420826 622454
rect 421062 622218 421146 622454
rect 421382 622218 421414 622454
rect 420794 622134 421414 622218
rect 420794 621898 420826 622134
rect 421062 621898 421146 622134
rect 421382 621898 421414 622134
rect 420794 582454 421414 621898
rect 420794 582218 420826 582454
rect 421062 582218 421146 582454
rect 421382 582218 421414 582454
rect 420794 582134 421414 582218
rect 420794 581898 420826 582134
rect 421062 581898 421146 582134
rect 421382 581898 421414 582134
rect 420794 542454 421414 581898
rect 420794 542218 420826 542454
rect 421062 542218 421146 542454
rect 421382 542218 421414 542454
rect 420794 542134 421414 542218
rect 420794 541898 420826 542134
rect 421062 541898 421146 542134
rect 421382 541898 421414 542134
rect 420794 502454 421414 541898
rect 420794 502218 420826 502454
rect 421062 502218 421146 502454
rect 421382 502218 421414 502454
rect 420794 502134 421414 502218
rect 420794 501898 420826 502134
rect 421062 501898 421146 502134
rect 421382 501898 421414 502134
rect 420794 462454 421414 501898
rect 420794 462218 420826 462454
rect 421062 462218 421146 462454
rect 421382 462218 421414 462454
rect 420794 462134 421414 462218
rect 420794 461898 420826 462134
rect 421062 461898 421146 462134
rect 421382 461898 421414 462134
rect 420794 422454 421414 461898
rect 420794 422218 420826 422454
rect 421062 422218 421146 422454
rect 421382 422218 421414 422454
rect 420794 422134 421414 422218
rect 420794 421898 420826 422134
rect 421062 421898 421146 422134
rect 421382 421898 421414 422134
rect 420794 382454 421414 421898
rect 420794 382218 420826 382454
rect 421062 382218 421146 382454
rect 421382 382218 421414 382454
rect 420794 382134 421414 382218
rect 420794 381898 420826 382134
rect 421062 381898 421146 382134
rect 421382 381898 421414 382134
rect 420794 342454 421414 381898
rect 420794 342218 420826 342454
rect 421062 342218 421146 342454
rect 421382 342218 421414 342454
rect 420794 342134 421414 342218
rect 420794 341898 420826 342134
rect 421062 341898 421146 342134
rect 421382 341898 421414 342134
rect 420794 302454 421414 341898
rect 420794 302218 420826 302454
rect 421062 302218 421146 302454
rect 421382 302218 421414 302454
rect 420794 302134 421414 302218
rect 420794 301898 420826 302134
rect 421062 301898 421146 302134
rect 421382 301898 421414 302134
rect 420794 262454 421414 301898
rect 420794 262218 420826 262454
rect 421062 262218 421146 262454
rect 421382 262218 421414 262454
rect 420794 262134 421414 262218
rect 420794 261898 420826 262134
rect 421062 261898 421146 262134
rect 421382 261898 421414 262134
rect 420794 222454 421414 261898
rect 420794 222218 420826 222454
rect 421062 222218 421146 222454
rect 421382 222218 421414 222454
rect 420794 222134 421414 222218
rect 420794 221898 420826 222134
rect 421062 221898 421146 222134
rect 421382 221898 421414 222134
rect 420794 182454 421414 221898
rect 420794 182218 420826 182454
rect 421062 182218 421146 182454
rect 421382 182218 421414 182454
rect 420794 182134 421414 182218
rect 420794 181898 420826 182134
rect 421062 181898 421146 182134
rect 421382 181898 421414 182134
rect 420794 142454 421414 181898
rect 420794 142218 420826 142454
rect 421062 142218 421146 142454
rect 421382 142218 421414 142454
rect 420794 142134 421414 142218
rect 420794 141898 420826 142134
rect 421062 141898 421146 142134
rect 421382 141898 421414 142134
rect 420794 102454 421414 141898
rect 420794 102218 420826 102454
rect 421062 102218 421146 102454
rect 421382 102218 421414 102454
rect 420794 102134 421414 102218
rect 420794 101898 420826 102134
rect 421062 101898 421146 102134
rect 421382 101898 421414 102134
rect 420794 62454 421414 101898
rect 420794 62218 420826 62454
rect 421062 62218 421146 62454
rect 421382 62218 421414 62454
rect 420794 62134 421414 62218
rect 420794 61898 420826 62134
rect 421062 61898 421146 62134
rect 421382 61898 421414 62134
rect 420794 22454 421414 61898
rect 420794 22218 420826 22454
rect 421062 22218 421146 22454
rect 421382 22218 421414 22454
rect 420794 22134 421414 22218
rect 420794 21898 420826 22134
rect 421062 21898 421146 22134
rect 421382 21898 421414 22134
rect 420794 -1306 421414 21898
rect 420794 -1542 420826 -1306
rect 421062 -1542 421146 -1306
rect 421382 -1542 421414 -1306
rect 420794 -1626 421414 -1542
rect 420794 -1862 420826 -1626
rect 421062 -1862 421146 -1626
rect 421382 -1862 421414 -1626
rect 420794 -1894 421414 -1862
rect 424514 666174 425134 707162
rect 424514 665938 424546 666174
rect 424782 665938 424866 666174
rect 425102 665938 425134 666174
rect 424514 665854 425134 665938
rect 424514 665618 424546 665854
rect 424782 665618 424866 665854
rect 425102 665618 425134 665854
rect 424514 626174 425134 665618
rect 424514 625938 424546 626174
rect 424782 625938 424866 626174
rect 425102 625938 425134 626174
rect 424514 625854 425134 625938
rect 424514 625618 424546 625854
rect 424782 625618 424866 625854
rect 425102 625618 425134 625854
rect 424514 586174 425134 625618
rect 424514 585938 424546 586174
rect 424782 585938 424866 586174
rect 425102 585938 425134 586174
rect 424514 585854 425134 585938
rect 424514 585618 424546 585854
rect 424782 585618 424866 585854
rect 425102 585618 425134 585854
rect 424514 546174 425134 585618
rect 424514 545938 424546 546174
rect 424782 545938 424866 546174
rect 425102 545938 425134 546174
rect 424514 545854 425134 545938
rect 424514 545618 424546 545854
rect 424782 545618 424866 545854
rect 425102 545618 425134 545854
rect 424514 506174 425134 545618
rect 424514 505938 424546 506174
rect 424782 505938 424866 506174
rect 425102 505938 425134 506174
rect 424514 505854 425134 505938
rect 424514 505618 424546 505854
rect 424782 505618 424866 505854
rect 425102 505618 425134 505854
rect 424514 466174 425134 505618
rect 424514 465938 424546 466174
rect 424782 465938 424866 466174
rect 425102 465938 425134 466174
rect 424514 465854 425134 465938
rect 424514 465618 424546 465854
rect 424782 465618 424866 465854
rect 425102 465618 425134 465854
rect 424514 426174 425134 465618
rect 424514 425938 424546 426174
rect 424782 425938 424866 426174
rect 425102 425938 425134 426174
rect 424514 425854 425134 425938
rect 424514 425618 424546 425854
rect 424782 425618 424866 425854
rect 425102 425618 425134 425854
rect 424514 386174 425134 425618
rect 424514 385938 424546 386174
rect 424782 385938 424866 386174
rect 425102 385938 425134 386174
rect 424514 385854 425134 385938
rect 424514 385618 424546 385854
rect 424782 385618 424866 385854
rect 425102 385618 425134 385854
rect 424514 346174 425134 385618
rect 424514 345938 424546 346174
rect 424782 345938 424866 346174
rect 425102 345938 425134 346174
rect 424514 345854 425134 345938
rect 424514 345618 424546 345854
rect 424782 345618 424866 345854
rect 425102 345618 425134 345854
rect 424514 306174 425134 345618
rect 424514 305938 424546 306174
rect 424782 305938 424866 306174
rect 425102 305938 425134 306174
rect 424514 305854 425134 305938
rect 424514 305618 424546 305854
rect 424782 305618 424866 305854
rect 425102 305618 425134 305854
rect 424514 266174 425134 305618
rect 424514 265938 424546 266174
rect 424782 265938 424866 266174
rect 425102 265938 425134 266174
rect 424514 265854 425134 265938
rect 424514 265618 424546 265854
rect 424782 265618 424866 265854
rect 425102 265618 425134 265854
rect 424514 226174 425134 265618
rect 424514 225938 424546 226174
rect 424782 225938 424866 226174
rect 425102 225938 425134 226174
rect 424514 225854 425134 225938
rect 424514 225618 424546 225854
rect 424782 225618 424866 225854
rect 425102 225618 425134 225854
rect 424514 186174 425134 225618
rect 424514 185938 424546 186174
rect 424782 185938 424866 186174
rect 425102 185938 425134 186174
rect 424514 185854 425134 185938
rect 424514 185618 424546 185854
rect 424782 185618 424866 185854
rect 425102 185618 425134 185854
rect 424514 146174 425134 185618
rect 424514 145938 424546 146174
rect 424782 145938 424866 146174
rect 425102 145938 425134 146174
rect 424514 145854 425134 145938
rect 424514 145618 424546 145854
rect 424782 145618 424866 145854
rect 425102 145618 425134 145854
rect 424514 106174 425134 145618
rect 424514 105938 424546 106174
rect 424782 105938 424866 106174
rect 425102 105938 425134 106174
rect 424514 105854 425134 105938
rect 424514 105618 424546 105854
rect 424782 105618 424866 105854
rect 425102 105618 425134 105854
rect 424514 66174 425134 105618
rect 424514 65938 424546 66174
rect 424782 65938 424866 66174
rect 425102 65938 425134 66174
rect 424514 65854 425134 65938
rect 424514 65618 424546 65854
rect 424782 65618 424866 65854
rect 425102 65618 425134 65854
rect 424514 26174 425134 65618
rect 424514 25938 424546 26174
rect 424782 25938 424866 26174
rect 425102 25938 425134 26174
rect 424514 25854 425134 25938
rect 424514 25618 424546 25854
rect 424782 25618 424866 25854
rect 425102 25618 425134 25854
rect 424514 -3226 425134 25618
rect 424514 -3462 424546 -3226
rect 424782 -3462 424866 -3226
rect 425102 -3462 425134 -3226
rect 424514 -3546 425134 -3462
rect 424514 -3782 424546 -3546
rect 424782 -3782 424866 -3546
rect 425102 -3782 425134 -3546
rect 424514 -3814 425134 -3782
rect 428234 669894 428854 709082
rect 428234 669658 428266 669894
rect 428502 669658 428586 669894
rect 428822 669658 428854 669894
rect 428234 669574 428854 669658
rect 428234 669338 428266 669574
rect 428502 669338 428586 669574
rect 428822 669338 428854 669574
rect 428234 629894 428854 669338
rect 428234 629658 428266 629894
rect 428502 629658 428586 629894
rect 428822 629658 428854 629894
rect 428234 629574 428854 629658
rect 428234 629338 428266 629574
rect 428502 629338 428586 629574
rect 428822 629338 428854 629574
rect 428234 589894 428854 629338
rect 428234 589658 428266 589894
rect 428502 589658 428586 589894
rect 428822 589658 428854 589894
rect 428234 589574 428854 589658
rect 428234 589338 428266 589574
rect 428502 589338 428586 589574
rect 428822 589338 428854 589574
rect 428234 549894 428854 589338
rect 428234 549658 428266 549894
rect 428502 549658 428586 549894
rect 428822 549658 428854 549894
rect 428234 549574 428854 549658
rect 428234 549338 428266 549574
rect 428502 549338 428586 549574
rect 428822 549338 428854 549574
rect 428234 509894 428854 549338
rect 428234 509658 428266 509894
rect 428502 509658 428586 509894
rect 428822 509658 428854 509894
rect 428234 509574 428854 509658
rect 428234 509338 428266 509574
rect 428502 509338 428586 509574
rect 428822 509338 428854 509574
rect 428234 469894 428854 509338
rect 428234 469658 428266 469894
rect 428502 469658 428586 469894
rect 428822 469658 428854 469894
rect 428234 469574 428854 469658
rect 428234 469338 428266 469574
rect 428502 469338 428586 469574
rect 428822 469338 428854 469574
rect 428234 429894 428854 469338
rect 428234 429658 428266 429894
rect 428502 429658 428586 429894
rect 428822 429658 428854 429894
rect 428234 429574 428854 429658
rect 428234 429338 428266 429574
rect 428502 429338 428586 429574
rect 428822 429338 428854 429574
rect 428234 389894 428854 429338
rect 428234 389658 428266 389894
rect 428502 389658 428586 389894
rect 428822 389658 428854 389894
rect 428234 389574 428854 389658
rect 428234 389338 428266 389574
rect 428502 389338 428586 389574
rect 428822 389338 428854 389574
rect 428234 349894 428854 389338
rect 428234 349658 428266 349894
rect 428502 349658 428586 349894
rect 428822 349658 428854 349894
rect 428234 349574 428854 349658
rect 428234 349338 428266 349574
rect 428502 349338 428586 349574
rect 428822 349338 428854 349574
rect 428234 309894 428854 349338
rect 428234 309658 428266 309894
rect 428502 309658 428586 309894
rect 428822 309658 428854 309894
rect 428234 309574 428854 309658
rect 428234 309338 428266 309574
rect 428502 309338 428586 309574
rect 428822 309338 428854 309574
rect 428234 269894 428854 309338
rect 428234 269658 428266 269894
rect 428502 269658 428586 269894
rect 428822 269658 428854 269894
rect 428234 269574 428854 269658
rect 428234 269338 428266 269574
rect 428502 269338 428586 269574
rect 428822 269338 428854 269574
rect 428234 229894 428854 269338
rect 428234 229658 428266 229894
rect 428502 229658 428586 229894
rect 428822 229658 428854 229894
rect 428234 229574 428854 229658
rect 428234 229338 428266 229574
rect 428502 229338 428586 229574
rect 428822 229338 428854 229574
rect 428234 189894 428854 229338
rect 428234 189658 428266 189894
rect 428502 189658 428586 189894
rect 428822 189658 428854 189894
rect 428234 189574 428854 189658
rect 428234 189338 428266 189574
rect 428502 189338 428586 189574
rect 428822 189338 428854 189574
rect 428234 149894 428854 189338
rect 428234 149658 428266 149894
rect 428502 149658 428586 149894
rect 428822 149658 428854 149894
rect 428234 149574 428854 149658
rect 428234 149338 428266 149574
rect 428502 149338 428586 149574
rect 428822 149338 428854 149574
rect 428234 109894 428854 149338
rect 428234 109658 428266 109894
rect 428502 109658 428586 109894
rect 428822 109658 428854 109894
rect 428234 109574 428854 109658
rect 428234 109338 428266 109574
rect 428502 109338 428586 109574
rect 428822 109338 428854 109574
rect 428234 69894 428854 109338
rect 428234 69658 428266 69894
rect 428502 69658 428586 69894
rect 428822 69658 428854 69894
rect 428234 69574 428854 69658
rect 428234 69338 428266 69574
rect 428502 69338 428586 69574
rect 428822 69338 428854 69574
rect 428234 29894 428854 69338
rect 428234 29658 428266 29894
rect 428502 29658 428586 29894
rect 428822 29658 428854 29894
rect 428234 29574 428854 29658
rect 428234 29338 428266 29574
rect 428502 29338 428586 29574
rect 428822 29338 428854 29574
rect 428234 -5146 428854 29338
rect 428234 -5382 428266 -5146
rect 428502 -5382 428586 -5146
rect 428822 -5382 428854 -5146
rect 428234 -5466 428854 -5382
rect 428234 -5702 428266 -5466
rect 428502 -5702 428586 -5466
rect 428822 -5702 428854 -5466
rect 428234 -5734 428854 -5702
rect 431954 673614 432574 711002
rect 451954 710598 452574 711590
rect 451954 710362 451986 710598
rect 452222 710362 452306 710598
rect 452542 710362 452574 710598
rect 451954 710278 452574 710362
rect 451954 710042 451986 710278
rect 452222 710042 452306 710278
rect 452542 710042 452574 710278
rect 448234 708678 448854 709670
rect 448234 708442 448266 708678
rect 448502 708442 448586 708678
rect 448822 708442 448854 708678
rect 448234 708358 448854 708442
rect 448234 708122 448266 708358
rect 448502 708122 448586 708358
rect 448822 708122 448854 708358
rect 444514 706758 445134 707750
rect 444514 706522 444546 706758
rect 444782 706522 444866 706758
rect 445102 706522 445134 706758
rect 444514 706438 445134 706522
rect 444514 706202 444546 706438
rect 444782 706202 444866 706438
rect 445102 706202 445134 706438
rect 431954 673378 431986 673614
rect 432222 673378 432306 673614
rect 432542 673378 432574 673614
rect 431954 673294 432574 673378
rect 431954 673058 431986 673294
rect 432222 673058 432306 673294
rect 432542 673058 432574 673294
rect 431954 633614 432574 673058
rect 431954 633378 431986 633614
rect 432222 633378 432306 633614
rect 432542 633378 432574 633614
rect 431954 633294 432574 633378
rect 431954 633058 431986 633294
rect 432222 633058 432306 633294
rect 432542 633058 432574 633294
rect 431954 593614 432574 633058
rect 431954 593378 431986 593614
rect 432222 593378 432306 593614
rect 432542 593378 432574 593614
rect 431954 593294 432574 593378
rect 431954 593058 431986 593294
rect 432222 593058 432306 593294
rect 432542 593058 432574 593294
rect 431954 553614 432574 593058
rect 431954 553378 431986 553614
rect 432222 553378 432306 553614
rect 432542 553378 432574 553614
rect 431954 553294 432574 553378
rect 431954 553058 431986 553294
rect 432222 553058 432306 553294
rect 432542 553058 432574 553294
rect 431954 513614 432574 553058
rect 431954 513378 431986 513614
rect 432222 513378 432306 513614
rect 432542 513378 432574 513614
rect 431954 513294 432574 513378
rect 431954 513058 431986 513294
rect 432222 513058 432306 513294
rect 432542 513058 432574 513294
rect 431954 473614 432574 513058
rect 431954 473378 431986 473614
rect 432222 473378 432306 473614
rect 432542 473378 432574 473614
rect 431954 473294 432574 473378
rect 431954 473058 431986 473294
rect 432222 473058 432306 473294
rect 432542 473058 432574 473294
rect 431954 433614 432574 473058
rect 431954 433378 431986 433614
rect 432222 433378 432306 433614
rect 432542 433378 432574 433614
rect 431954 433294 432574 433378
rect 431954 433058 431986 433294
rect 432222 433058 432306 433294
rect 432542 433058 432574 433294
rect 431954 393614 432574 433058
rect 431954 393378 431986 393614
rect 432222 393378 432306 393614
rect 432542 393378 432574 393614
rect 431954 393294 432574 393378
rect 431954 393058 431986 393294
rect 432222 393058 432306 393294
rect 432542 393058 432574 393294
rect 431954 353614 432574 393058
rect 431954 353378 431986 353614
rect 432222 353378 432306 353614
rect 432542 353378 432574 353614
rect 431954 353294 432574 353378
rect 431954 353058 431986 353294
rect 432222 353058 432306 353294
rect 432542 353058 432574 353294
rect 431954 313614 432574 353058
rect 431954 313378 431986 313614
rect 432222 313378 432306 313614
rect 432542 313378 432574 313614
rect 431954 313294 432574 313378
rect 431954 313058 431986 313294
rect 432222 313058 432306 313294
rect 432542 313058 432574 313294
rect 431954 273614 432574 313058
rect 431954 273378 431986 273614
rect 432222 273378 432306 273614
rect 432542 273378 432574 273614
rect 431954 273294 432574 273378
rect 431954 273058 431986 273294
rect 432222 273058 432306 273294
rect 432542 273058 432574 273294
rect 431954 233614 432574 273058
rect 431954 233378 431986 233614
rect 432222 233378 432306 233614
rect 432542 233378 432574 233614
rect 431954 233294 432574 233378
rect 431954 233058 431986 233294
rect 432222 233058 432306 233294
rect 432542 233058 432574 233294
rect 431954 193614 432574 233058
rect 431954 193378 431986 193614
rect 432222 193378 432306 193614
rect 432542 193378 432574 193614
rect 431954 193294 432574 193378
rect 431954 193058 431986 193294
rect 432222 193058 432306 193294
rect 432542 193058 432574 193294
rect 431954 153614 432574 193058
rect 431954 153378 431986 153614
rect 432222 153378 432306 153614
rect 432542 153378 432574 153614
rect 431954 153294 432574 153378
rect 431954 153058 431986 153294
rect 432222 153058 432306 153294
rect 432542 153058 432574 153294
rect 431954 113614 432574 153058
rect 431954 113378 431986 113614
rect 432222 113378 432306 113614
rect 432542 113378 432574 113614
rect 431954 113294 432574 113378
rect 431954 113058 431986 113294
rect 432222 113058 432306 113294
rect 432542 113058 432574 113294
rect 431954 73614 432574 113058
rect 431954 73378 431986 73614
rect 432222 73378 432306 73614
rect 432542 73378 432574 73614
rect 431954 73294 432574 73378
rect 431954 73058 431986 73294
rect 432222 73058 432306 73294
rect 432542 73058 432574 73294
rect 431954 33614 432574 73058
rect 431954 33378 431986 33614
rect 432222 33378 432306 33614
rect 432542 33378 432574 33614
rect 431954 33294 432574 33378
rect 431954 33058 431986 33294
rect 432222 33058 432306 33294
rect 432542 33058 432574 33294
rect 411954 -6342 411986 -6106
rect 412222 -6342 412306 -6106
rect 412542 -6342 412574 -6106
rect 411954 -6426 412574 -6342
rect 411954 -6662 411986 -6426
rect 412222 -6662 412306 -6426
rect 412542 -6662 412574 -6426
rect 411954 -7654 412574 -6662
rect 431954 -7066 432574 33058
rect 440794 704838 441414 705830
rect 440794 704602 440826 704838
rect 441062 704602 441146 704838
rect 441382 704602 441414 704838
rect 440794 704518 441414 704602
rect 440794 704282 440826 704518
rect 441062 704282 441146 704518
rect 441382 704282 441414 704518
rect 440794 682454 441414 704282
rect 440794 682218 440826 682454
rect 441062 682218 441146 682454
rect 441382 682218 441414 682454
rect 440794 682134 441414 682218
rect 440794 681898 440826 682134
rect 441062 681898 441146 682134
rect 441382 681898 441414 682134
rect 440794 642454 441414 681898
rect 440794 642218 440826 642454
rect 441062 642218 441146 642454
rect 441382 642218 441414 642454
rect 440794 642134 441414 642218
rect 440794 641898 440826 642134
rect 441062 641898 441146 642134
rect 441382 641898 441414 642134
rect 440794 602454 441414 641898
rect 440794 602218 440826 602454
rect 441062 602218 441146 602454
rect 441382 602218 441414 602454
rect 440794 602134 441414 602218
rect 440794 601898 440826 602134
rect 441062 601898 441146 602134
rect 441382 601898 441414 602134
rect 440794 562454 441414 601898
rect 440794 562218 440826 562454
rect 441062 562218 441146 562454
rect 441382 562218 441414 562454
rect 440794 562134 441414 562218
rect 440794 561898 440826 562134
rect 441062 561898 441146 562134
rect 441382 561898 441414 562134
rect 440794 522454 441414 561898
rect 440794 522218 440826 522454
rect 441062 522218 441146 522454
rect 441382 522218 441414 522454
rect 440794 522134 441414 522218
rect 440794 521898 440826 522134
rect 441062 521898 441146 522134
rect 441382 521898 441414 522134
rect 440794 482454 441414 521898
rect 440794 482218 440826 482454
rect 441062 482218 441146 482454
rect 441382 482218 441414 482454
rect 440794 482134 441414 482218
rect 440794 481898 440826 482134
rect 441062 481898 441146 482134
rect 441382 481898 441414 482134
rect 440794 442454 441414 481898
rect 440794 442218 440826 442454
rect 441062 442218 441146 442454
rect 441382 442218 441414 442454
rect 440794 442134 441414 442218
rect 440794 441898 440826 442134
rect 441062 441898 441146 442134
rect 441382 441898 441414 442134
rect 440794 402454 441414 441898
rect 440794 402218 440826 402454
rect 441062 402218 441146 402454
rect 441382 402218 441414 402454
rect 440794 402134 441414 402218
rect 440794 401898 440826 402134
rect 441062 401898 441146 402134
rect 441382 401898 441414 402134
rect 440794 362454 441414 401898
rect 440794 362218 440826 362454
rect 441062 362218 441146 362454
rect 441382 362218 441414 362454
rect 440794 362134 441414 362218
rect 440794 361898 440826 362134
rect 441062 361898 441146 362134
rect 441382 361898 441414 362134
rect 440794 322454 441414 361898
rect 440794 322218 440826 322454
rect 441062 322218 441146 322454
rect 441382 322218 441414 322454
rect 440794 322134 441414 322218
rect 440794 321898 440826 322134
rect 441062 321898 441146 322134
rect 441382 321898 441414 322134
rect 440794 282454 441414 321898
rect 440794 282218 440826 282454
rect 441062 282218 441146 282454
rect 441382 282218 441414 282454
rect 440794 282134 441414 282218
rect 440794 281898 440826 282134
rect 441062 281898 441146 282134
rect 441382 281898 441414 282134
rect 440794 242454 441414 281898
rect 440794 242218 440826 242454
rect 441062 242218 441146 242454
rect 441382 242218 441414 242454
rect 440794 242134 441414 242218
rect 440794 241898 440826 242134
rect 441062 241898 441146 242134
rect 441382 241898 441414 242134
rect 440794 202454 441414 241898
rect 440794 202218 440826 202454
rect 441062 202218 441146 202454
rect 441382 202218 441414 202454
rect 440794 202134 441414 202218
rect 440794 201898 440826 202134
rect 441062 201898 441146 202134
rect 441382 201898 441414 202134
rect 440794 162454 441414 201898
rect 440794 162218 440826 162454
rect 441062 162218 441146 162454
rect 441382 162218 441414 162454
rect 440794 162134 441414 162218
rect 440794 161898 440826 162134
rect 441062 161898 441146 162134
rect 441382 161898 441414 162134
rect 440794 122454 441414 161898
rect 440794 122218 440826 122454
rect 441062 122218 441146 122454
rect 441382 122218 441414 122454
rect 440794 122134 441414 122218
rect 440794 121898 440826 122134
rect 441062 121898 441146 122134
rect 441382 121898 441414 122134
rect 440794 82454 441414 121898
rect 440794 82218 440826 82454
rect 441062 82218 441146 82454
rect 441382 82218 441414 82454
rect 440794 82134 441414 82218
rect 440794 81898 440826 82134
rect 441062 81898 441146 82134
rect 441382 81898 441414 82134
rect 440794 42454 441414 81898
rect 440794 42218 440826 42454
rect 441062 42218 441146 42454
rect 441382 42218 441414 42454
rect 440794 42134 441414 42218
rect 440794 41898 440826 42134
rect 441062 41898 441146 42134
rect 441382 41898 441414 42134
rect 440794 2454 441414 41898
rect 440794 2218 440826 2454
rect 441062 2218 441146 2454
rect 441382 2218 441414 2454
rect 440794 2134 441414 2218
rect 440794 1898 440826 2134
rect 441062 1898 441146 2134
rect 441382 1898 441414 2134
rect 440794 -346 441414 1898
rect 440794 -582 440826 -346
rect 441062 -582 441146 -346
rect 441382 -582 441414 -346
rect 440794 -666 441414 -582
rect 440794 -902 440826 -666
rect 441062 -902 441146 -666
rect 441382 -902 441414 -666
rect 440794 -1894 441414 -902
rect 444514 686174 445134 706202
rect 444514 685938 444546 686174
rect 444782 685938 444866 686174
rect 445102 685938 445134 686174
rect 444514 685854 445134 685938
rect 444514 685618 444546 685854
rect 444782 685618 444866 685854
rect 445102 685618 445134 685854
rect 444514 646174 445134 685618
rect 444514 645938 444546 646174
rect 444782 645938 444866 646174
rect 445102 645938 445134 646174
rect 444514 645854 445134 645938
rect 444514 645618 444546 645854
rect 444782 645618 444866 645854
rect 445102 645618 445134 645854
rect 444514 606174 445134 645618
rect 444514 605938 444546 606174
rect 444782 605938 444866 606174
rect 445102 605938 445134 606174
rect 444514 605854 445134 605938
rect 444514 605618 444546 605854
rect 444782 605618 444866 605854
rect 445102 605618 445134 605854
rect 444514 566174 445134 605618
rect 444514 565938 444546 566174
rect 444782 565938 444866 566174
rect 445102 565938 445134 566174
rect 444514 565854 445134 565938
rect 444514 565618 444546 565854
rect 444782 565618 444866 565854
rect 445102 565618 445134 565854
rect 444514 526174 445134 565618
rect 444514 525938 444546 526174
rect 444782 525938 444866 526174
rect 445102 525938 445134 526174
rect 444514 525854 445134 525938
rect 444514 525618 444546 525854
rect 444782 525618 444866 525854
rect 445102 525618 445134 525854
rect 444514 486174 445134 525618
rect 444514 485938 444546 486174
rect 444782 485938 444866 486174
rect 445102 485938 445134 486174
rect 444514 485854 445134 485938
rect 444514 485618 444546 485854
rect 444782 485618 444866 485854
rect 445102 485618 445134 485854
rect 444514 446174 445134 485618
rect 444514 445938 444546 446174
rect 444782 445938 444866 446174
rect 445102 445938 445134 446174
rect 444514 445854 445134 445938
rect 444514 445618 444546 445854
rect 444782 445618 444866 445854
rect 445102 445618 445134 445854
rect 444514 406174 445134 445618
rect 444514 405938 444546 406174
rect 444782 405938 444866 406174
rect 445102 405938 445134 406174
rect 444514 405854 445134 405938
rect 444514 405618 444546 405854
rect 444782 405618 444866 405854
rect 445102 405618 445134 405854
rect 444514 366174 445134 405618
rect 444514 365938 444546 366174
rect 444782 365938 444866 366174
rect 445102 365938 445134 366174
rect 444514 365854 445134 365938
rect 444514 365618 444546 365854
rect 444782 365618 444866 365854
rect 445102 365618 445134 365854
rect 444514 326174 445134 365618
rect 444514 325938 444546 326174
rect 444782 325938 444866 326174
rect 445102 325938 445134 326174
rect 444514 325854 445134 325938
rect 444514 325618 444546 325854
rect 444782 325618 444866 325854
rect 445102 325618 445134 325854
rect 444514 286174 445134 325618
rect 444514 285938 444546 286174
rect 444782 285938 444866 286174
rect 445102 285938 445134 286174
rect 444514 285854 445134 285938
rect 444514 285618 444546 285854
rect 444782 285618 444866 285854
rect 445102 285618 445134 285854
rect 444514 246174 445134 285618
rect 444514 245938 444546 246174
rect 444782 245938 444866 246174
rect 445102 245938 445134 246174
rect 444514 245854 445134 245938
rect 444514 245618 444546 245854
rect 444782 245618 444866 245854
rect 445102 245618 445134 245854
rect 444514 206174 445134 245618
rect 444514 205938 444546 206174
rect 444782 205938 444866 206174
rect 445102 205938 445134 206174
rect 444514 205854 445134 205938
rect 444514 205618 444546 205854
rect 444782 205618 444866 205854
rect 445102 205618 445134 205854
rect 444514 166174 445134 205618
rect 444514 165938 444546 166174
rect 444782 165938 444866 166174
rect 445102 165938 445134 166174
rect 444514 165854 445134 165938
rect 444514 165618 444546 165854
rect 444782 165618 444866 165854
rect 445102 165618 445134 165854
rect 444514 126174 445134 165618
rect 444514 125938 444546 126174
rect 444782 125938 444866 126174
rect 445102 125938 445134 126174
rect 444514 125854 445134 125938
rect 444514 125618 444546 125854
rect 444782 125618 444866 125854
rect 445102 125618 445134 125854
rect 444514 86174 445134 125618
rect 444514 85938 444546 86174
rect 444782 85938 444866 86174
rect 445102 85938 445134 86174
rect 444514 85854 445134 85938
rect 444514 85618 444546 85854
rect 444782 85618 444866 85854
rect 445102 85618 445134 85854
rect 444514 46174 445134 85618
rect 444514 45938 444546 46174
rect 444782 45938 444866 46174
rect 445102 45938 445134 46174
rect 444514 45854 445134 45938
rect 444514 45618 444546 45854
rect 444782 45618 444866 45854
rect 445102 45618 445134 45854
rect 444514 6174 445134 45618
rect 444514 5938 444546 6174
rect 444782 5938 444866 6174
rect 445102 5938 445134 6174
rect 444514 5854 445134 5938
rect 444514 5618 444546 5854
rect 444782 5618 444866 5854
rect 445102 5618 445134 5854
rect 444514 -2266 445134 5618
rect 444514 -2502 444546 -2266
rect 444782 -2502 444866 -2266
rect 445102 -2502 445134 -2266
rect 444514 -2586 445134 -2502
rect 444514 -2822 444546 -2586
rect 444782 -2822 444866 -2586
rect 445102 -2822 445134 -2586
rect 444514 -3814 445134 -2822
rect 448234 689894 448854 708122
rect 448234 689658 448266 689894
rect 448502 689658 448586 689894
rect 448822 689658 448854 689894
rect 448234 689574 448854 689658
rect 448234 689338 448266 689574
rect 448502 689338 448586 689574
rect 448822 689338 448854 689574
rect 448234 649894 448854 689338
rect 448234 649658 448266 649894
rect 448502 649658 448586 649894
rect 448822 649658 448854 649894
rect 448234 649574 448854 649658
rect 448234 649338 448266 649574
rect 448502 649338 448586 649574
rect 448822 649338 448854 649574
rect 448234 609894 448854 649338
rect 448234 609658 448266 609894
rect 448502 609658 448586 609894
rect 448822 609658 448854 609894
rect 448234 609574 448854 609658
rect 448234 609338 448266 609574
rect 448502 609338 448586 609574
rect 448822 609338 448854 609574
rect 448234 569894 448854 609338
rect 448234 569658 448266 569894
rect 448502 569658 448586 569894
rect 448822 569658 448854 569894
rect 448234 569574 448854 569658
rect 448234 569338 448266 569574
rect 448502 569338 448586 569574
rect 448822 569338 448854 569574
rect 448234 529894 448854 569338
rect 448234 529658 448266 529894
rect 448502 529658 448586 529894
rect 448822 529658 448854 529894
rect 448234 529574 448854 529658
rect 448234 529338 448266 529574
rect 448502 529338 448586 529574
rect 448822 529338 448854 529574
rect 448234 489894 448854 529338
rect 448234 489658 448266 489894
rect 448502 489658 448586 489894
rect 448822 489658 448854 489894
rect 448234 489574 448854 489658
rect 448234 489338 448266 489574
rect 448502 489338 448586 489574
rect 448822 489338 448854 489574
rect 448234 449894 448854 489338
rect 448234 449658 448266 449894
rect 448502 449658 448586 449894
rect 448822 449658 448854 449894
rect 448234 449574 448854 449658
rect 448234 449338 448266 449574
rect 448502 449338 448586 449574
rect 448822 449338 448854 449574
rect 448234 409894 448854 449338
rect 448234 409658 448266 409894
rect 448502 409658 448586 409894
rect 448822 409658 448854 409894
rect 448234 409574 448854 409658
rect 448234 409338 448266 409574
rect 448502 409338 448586 409574
rect 448822 409338 448854 409574
rect 448234 369894 448854 409338
rect 448234 369658 448266 369894
rect 448502 369658 448586 369894
rect 448822 369658 448854 369894
rect 448234 369574 448854 369658
rect 448234 369338 448266 369574
rect 448502 369338 448586 369574
rect 448822 369338 448854 369574
rect 448234 329894 448854 369338
rect 448234 329658 448266 329894
rect 448502 329658 448586 329894
rect 448822 329658 448854 329894
rect 448234 329574 448854 329658
rect 448234 329338 448266 329574
rect 448502 329338 448586 329574
rect 448822 329338 448854 329574
rect 448234 289894 448854 329338
rect 448234 289658 448266 289894
rect 448502 289658 448586 289894
rect 448822 289658 448854 289894
rect 448234 289574 448854 289658
rect 448234 289338 448266 289574
rect 448502 289338 448586 289574
rect 448822 289338 448854 289574
rect 448234 249894 448854 289338
rect 448234 249658 448266 249894
rect 448502 249658 448586 249894
rect 448822 249658 448854 249894
rect 448234 249574 448854 249658
rect 448234 249338 448266 249574
rect 448502 249338 448586 249574
rect 448822 249338 448854 249574
rect 448234 209894 448854 249338
rect 448234 209658 448266 209894
rect 448502 209658 448586 209894
rect 448822 209658 448854 209894
rect 448234 209574 448854 209658
rect 448234 209338 448266 209574
rect 448502 209338 448586 209574
rect 448822 209338 448854 209574
rect 448234 169894 448854 209338
rect 448234 169658 448266 169894
rect 448502 169658 448586 169894
rect 448822 169658 448854 169894
rect 448234 169574 448854 169658
rect 448234 169338 448266 169574
rect 448502 169338 448586 169574
rect 448822 169338 448854 169574
rect 448234 129894 448854 169338
rect 448234 129658 448266 129894
rect 448502 129658 448586 129894
rect 448822 129658 448854 129894
rect 448234 129574 448854 129658
rect 448234 129338 448266 129574
rect 448502 129338 448586 129574
rect 448822 129338 448854 129574
rect 448234 89894 448854 129338
rect 448234 89658 448266 89894
rect 448502 89658 448586 89894
rect 448822 89658 448854 89894
rect 448234 89574 448854 89658
rect 448234 89338 448266 89574
rect 448502 89338 448586 89574
rect 448822 89338 448854 89574
rect 448234 49894 448854 89338
rect 448234 49658 448266 49894
rect 448502 49658 448586 49894
rect 448822 49658 448854 49894
rect 448234 49574 448854 49658
rect 448234 49338 448266 49574
rect 448502 49338 448586 49574
rect 448822 49338 448854 49574
rect 448234 9894 448854 49338
rect 448234 9658 448266 9894
rect 448502 9658 448586 9894
rect 448822 9658 448854 9894
rect 448234 9574 448854 9658
rect 448234 9338 448266 9574
rect 448502 9338 448586 9574
rect 448822 9338 448854 9574
rect 448234 -4186 448854 9338
rect 448234 -4422 448266 -4186
rect 448502 -4422 448586 -4186
rect 448822 -4422 448854 -4186
rect 448234 -4506 448854 -4422
rect 448234 -4742 448266 -4506
rect 448502 -4742 448586 -4506
rect 448822 -4742 448854 -4506
rect 448234 -5734 448854 -4742
rect 451954 693614 452574 710042
rect 471954 711558 472574 711590
rect 471954 711322 471986 711558
rect 472222 711322 472306 711558
rect 472542 711322 472574 711558
rect 471954 711238 472574 711322
rect 471954 711002 471986 711238
rect 472222 711002 472306 711238
rect 472542 711002 472574 711238
rect 468234 709638 468854 709670
rect 468234 709402 468266 709638
rect 468502 709402 468586 709638
rect 468822 709402 468854 709638
rect 468234 709318 468854 709402
rect 468234 709082 468266 709318
rect 468502 709082 468586 709318
rect 468822 709082 468854 709318
rect 464514 707718 465134 707750
rect 464514 707482 464546 707718
rect 464782 707482 464866 707718
rect 465102 707482 465134 707718
rect 464514 707398 465134 707482
rect 464514 707162 464546 707398
rect 464782 707162 464866 707398
rect 465102 707162 465134 707398
rect 451954 693378 451986 693614
rect 452222 693378 452306 693614
rect 452542 693378 452574 693614
rect 451954 693294 452574 693378
rect 451954 693058 451986 693294
rect 452222 693058 452306 693294
rect 452542 693058 452574 693294
rect 451954 653614 452574 693058
rect 451954 653378 451986 653614
rect 452222 653378 452306 653614
rect 452542 653378 452574 653614
rect 451954 653294 452574 653378
rect 451954 653058 451986 653294
rect 452222 653058 452306 653294
rect 452542 653058 452574 653294
rect 451954 613614 452574 653058
rect 451954 613378 451986 613614
rect 452222 613378 452306 613614
rect 452542 613378 452574 613614
rect 451954 613294 452574 613378
rect 451954 613058 451986 613294
rect 452222 613058 452306 613294
rect 452542 613058 452574 613294
rect 451954 573614 452574 613058
rect 451954 573378 451986 573614
rect 452222 573378 452306 573614
rect 452542 573378 452574 573614
rect 451954 573294 452574 573378
rect 451954 573058 451986 573294
rect 452222 573058 452306 573294
rect 452542 573058 452574 573294
rect 451954 533614 452574 573058
rect 451954 533378 451986 533614
rect 452222 533378 452306 533614
rect 452542 533378 452574 533614
rect 451954 533294 452574 533378
rect 451954 533058 451986 533294
rect 452222 533058 452306 533294
rect 452542 533058 452574 533294
rect 451954 493614 452574 533058
rect 451954 493378 451986 493614
rect 452222 493378 452306 493614
rect 452542 493378 452574 493614
rect 451954 493294 452574 493378
rect 451954 493058 451986 493294
rect 452222 493058 452306 493294
rect 452542 493058 452574 493294
rect 451954 453614 452574 493058
rect 451954 453378 451986 453614
rect 452222 453378 452306 453614
rect 452542 453378 452574 453614
rect 451954 453294 452574 453378
rect 451954 453058 451986 453294
rect 452222 453058 452306 453294
rect 452542 453058 452574 453294
rect 451954 413614 452574 453058
rect 451954 413378 451986 413614
rect 452222 413378 452306 413614
rect 452542 413378 452574 413614
rect 451954 413294 452574 413378
rect 451954 413058 451986 413294
rect 452222 413058 452306 413294
rect 452542 413058 452574 413294
rect 451954 373614 452574 413058
rect 451954 373378 451986 373614
rect 452222 373378 452306 373614
rect 452542 373378 452574 373614
rect 451954 373294 452574 373378
rect 451954 373058 451986 373294
rect 452222 373058 452306 373294
rect 452542 373058 452574 373294
rect 451954 333614 452574 373058
rect 451954 333378 451986 333614
rect 452222 333378 452306 333614
rect 452542 333378 452574 333614
rect 451954 333294 452574 333378
rect 451954 333058 451986 333294
rect 452222 333058 452306 333294
rect 452542 333058 452574 333294
rect 451954 293614 452574 333058
rect 451954 293378 451986 293614
rect 452222 293378 452306 293614
rect 452542 293378 452574 293614
rect 451954 293294 452574 293378
rect 451954 293058 451986 293294
rect 452222 293058 452306 293294
rect 452542 293058 452574 293294
rect 451954 253614 452574 293058
rect 451954 253378 451986 253614
rect 452222 253378 452306 253614
rect 452542 253378 452574 253614
rect 451954 253294 452574 253378
rect 451954 253058 451986 253294
rect 452222 253058 452306 253294
rect 452542 253058 452574 253294
rect 451954 213614 452574 253058
rect 451954 213378 451986 213614
rect 452222 213378 452306 213614
rect 452542 213378 452574 213614
rect 451954 213294 452574 213378
rect 451954 213058 451986 213294
rect 452222 213058 452306 213294
rect 452542 213058 452574 213294
rect 451954 173614 452574 213058
rect 451954 173378 451986 173614
rect 452222 173378 452306 173614
rect 452542 173378 452574 173614
rect 451954 173294 452574 173378
rect 451954 173058 451986 173294
rect 452222 173058 452306 173294
rect 452542 173058 452574 173294
rect 451954 133614 452574 173058
rect 451954 133378 451986 133614
rect 452222 133378 452306 133614
rect 452542 133378 452574 133614
rect 451954 133294 452574 133378
rect 451954 133058 451986 133294
rect 452222 133058 452306 133294
rect 452542 133058 452574 133294
rect 451954 93614 452574 133058
rect 451954 93378 451986 93614
rect 452222 93378 452306 93614
rect 452542 93378 452574 93614
rect 451954 93294 452574 93378
rect 451954 93058 451986 93294
rect 452222 93058 452306 93294
rect 452542 93058 452574 93294
rect 451954 53614 452574 93058
rect 451954 53378 451986 53614
rect 452222 53378 452306 53614
rect 452542 53378 452574 53614
rect 451954 53294 452574 53378
rect 451954 53058 451986 53294
rect 452222 53058 452306 53294
rect 452542 53058 452574 53294
rect 451954 13614 452574 53058
rect 451954 13378 451986 13614
rect 452222 13378 452306 13614
rect 452542 13378 452574 13614
rect 451954 13294 452574 13378
rect 451954 13058 451986 13294
rect 452222 13058 452306 13294
rect 452542 13058 452574 13294
rect 431954 -7302 431986 -7066
rect 432222 -7302 432306 -7066
rect 432542 -7302 432574 -7066
rect 431954 -7386 432574 -7302
rect 431954 -7622 431986 -7386
rect 432222 -7622 432306 -7386
rect 432542 -7622 432574 -7386
rect 431954 -7654 432574 -7622
rect 451954 -6106 452574 13058
rect 460794 705798 461414 705830
rect 460794 705562 460826 705798
rect 461062 705562 461146 705798
rect 461382 705562 461414 705798
rect 460794 705478 461414 705562
rect 460794 705242 460826 705478
rect 461062 705242 461146 705478
rect 461382 705242 461414 705478
rect 460794 662454 461414 705242
rect 460794 662218 460826 662454
rect 461062 662218 461146 662454
rect 461382 662218 461414 662454
rect 460794 662134 461414 662218
rect 460794 661898 460826 662134
rect 461062 661898 461146 662134
rect 461382 661898 461414 662134
rect 460794 622454 461414 661898
rect 460794 622218 460826 622454
rect 461062 622218 461146 622454
rect 461382 622218 461414 622454
rect 460794 622134 461414 622218
rect 460794 621898 460826 622134
rect 461062 621898 461146 622134
rect 461382 621898 461414 622134
rect 460794 582454 461414 621898
rect 460794 582218 460826 582454
rect 461062 582218 461146 582454
rect 461382 582218 461414 582454
rect 460794 582134 461414 582218
rect 460794 581898 460826 582134
rect 461062 581898 461146 582134
rect 461382 581898 461414 582134
rect 460794 542454 461414 581898
rect 460794 542218 460826 542454
rect 461062 542218 461146 542454
rect 461382 542218 461414 542454
rect 460794 542134 461414 542218
rect 460794 541898 460826 542134
rect 461062 541898 461146 542134
rect 461382 541898 461414 542134
rect 460794 502454 461414 541898
rect 460794 502218 460826 502454
rect 461062 502218 461146 502454
rect 461382 502218 461414 502454
rect 460794 502134 461414 502218
rect 460794 501898 460826 502134
rect 461062 501898 461146 502134
rect 461382 501898 461414 502134
rect 460794 462454 461414 501898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 422454 461414 461898
rect 460794 422218 460826 422454
rect 461062 422218 461146 422454
rect 461382 422218 461414 422454
rect 460794 422134 461414 422218
rect 460794 421898 460826 422134
rect 461062 421898 461146 422134
rect 461382 421898 461414 422134
rect 460794 382454 461414 421898
rect 460794 382218 460826 382454
rect 461062 382218 461146 382454
rect 461382 382218 461414 382454
rect 460794 382134 461414 382218
rect 460794 381898 460826 382134
rect 461062 381898 461146 382134
rect 461382 381898 461414 382134
rect 460794 342454 461414 381898
rect 460794 342218 460826 342454
rect 461062 342218 461146 342454
rect 461382 342218 461414 342454
rect 460794 342134 461414 342218
rect 460794 341898 460826 342134
rect 461062 341898 461146 342134
rect 461382 341898 461414 342134
rect 460794 302454 461414 341898
rect 460794 302218 460826 302454
rect 461062 302218 461146 302454
rect 461382 302218 461414 302454
rect 460794 302134 461414 302218
rect 460794 301898 460826 302134
rect 461062 301898 461146 302134
rect 461382 301898 461414 302134
rect 460794 262454 461414 301898
rect 460794 262218 460826 262454
rect 461062 262218 461146 262454
rect 461382 262218 461414 262454
rect 460794 262134 461414 262218
rect 460794 261898 460826 262134
rect 461062 261898 461146 262134
rect 461382 261898 461414 262134
rect 460794 222454 461414 261898
rect 460794 222218 460826 222454
rect 461062 222218 461146 222454
rect 461382 222218 461414 222454
rect 460794 222134 461414 222218
rect 460794 221898 460826 222134
rect 461062 221898 461146 222134
rect 461382 221898 461414 222134
rect 460794 182454 461414 221898
rect 460794 182218 460826 182454
rect 461062 182218 461146 182454
rect 461382 182218 461414 182454
rect 460794 182134 461414 182218
rect 460794 181898 460826 182134
rect 461062 181898 461146 182134
rect 461382 181898 461414 182134
rect 460794 142454 461414 181898
rect 460794 142218 460826 142454
rect 461062 142218 461146 142454
rect 461382 142218 461414 142454
rect 460794 142134 461414 142218
rect 460794 141898 460826 142134
rect 461062 141898 461146 142134
rect 461382 141898 461414 142134
rect 460794 102454 461414 141898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 62454 461414 101898
rect 460794 62218 460826 62454
rect 461062 62218 461146 62454
rect 461382 62218 461414 62454
rect 460794 62134 461414 62218
rect 460794 61898 460826 62134
rect 461062 61898 461146 62134
rect 461382 61898 461414 62134
rect 460794 22454 461414 61898
rect 460794 22218 460826 22454
rect 461062 22218 461146 22454
rect 461382 22218 461414 22454
rect 460794 22134 461414 22218
rect 460794 21898 460826 22134
rect 461062 21898 461146 22134
rect 461382 21898 461414 22134
rect 460794 -1306 461414 21898
rect 460794 -1542 460826 -1306
rect 461062 -1542 461146 -1306
rect 461382 -1542 461414 -1306
rect 460794 -1626 461414 -1542
rect 460794 -1862 460826 -1626
rect 461062 -1862 461146 -1626
rect 461382 -1862 461414 -1626
rect 460794 -1894 461414 -1862
rect 464514 666174 465134 707162
rect 464514 665938 464546 666174
rect 464782 665938 464866 666174
rect 465102 665938 465134 666174
rect 464514 665854 465134 665938
rect 464514 665618 464546 665854
rect 464782 665618 464866 665854
rect 465102 665618 465134 665854
rect 464514 626174 465134 665618
rect 464514 625938 464546 626174
rect 464782 625938 464866 626174
rect 465102 625938 465134 626174
rect 464514 625854 465134 625938
rect 464514 625618 464546 625854
rect 464782 625618 464866 625854
rect 465102 625618 465134 625854
rect 464514 586174 465134 625618
rect 464514 585938 464546 586174
rect 464782 585938 464866 586174
rect 465102 585938 465134 586174
rect 464514 585854 465134 585938
rect 464514 585618 464546 585854
rect 464782 585618 464866 585854
rect 465102 585618 465134 585854
rect 464514 546174 465134 585618
rect 464514 545938 464546 546174
rect 464782 545938 464866 546174
rect 465102 545938 465134 546174
rect 464514 545854 465134 545938
rect 464514 545618 464546 545854
rect 464782 545618 464866 545854
rect 465102 545618 465134 545854
rect 464514 506174 465134 545618
rect 464514 505938 464546 506174
rect 464782 505938 464866 506174
rect 465102 505938 465134 506174
rect 464514 505854 465134 505938
rect 464514 505618 464546 505854
rect 464782 505618 464866 505854
rect 465102 505618 465134 505854
rect 464514 466174 465134 505618
rect 464514 465938 464546 466174
rect 464782 465938 464866 466174
rect 465102 465938 465134 466174
rect 464514 465854 465134 465938
rect 464514 465618 464546 465854
rect 464782 465618 464866 465854
rect 465102 465618 465134 465854
rect 464514 426174 465134 465618
rect 464514 425938 464546 426174
rect 464782 425938 464866 426174
rect 465102 425938 465134 426174
rect 464514 425854 465134 425938
rect 464514 425618 464546 425854
rect 464782 425618 464866 425854
rect 465102 425618 465134 425854
rect 464514 386174 465134 425618
rect 464514 385938 464546 386174
rect 464782 385938 464866 386174
rect 465102 385938 465134 386174
rect 464514 385854 465134 385938
rect 464514 385618 464546 385854
rect 464782 385618 464866 385854
rect 465102 385618 465134 385854
rect 464514 346174 465134 385618
rect 464514 345938 464546 346174
rect 464782 345938 464866 346174
rect 465102 345938 465134 346174
rect 464514 345854 465134 345938
rect 464514 345618 464546 345854
rect 464782 345618 464866 345854
rect 465102 345618 465134 345854
rect 464514 306174 465134 345618
rect 464514 305938 464546 306174
rect 464782 305938 464866 306174
rect 465102 305938 465134 306174
rect 464514 305854 465134 305938
rect 464514 305618 464546 305854
rect 464782 305618 464866 305854
rect 465102 305618 465134 305854
rect 464514 266174 465134 305618
rect 464514 265938 464546 266174
rect 464782 265938 464866 266174
rect 465102 265938 465134 266174
rect 464514 265854 465134 265938
rect 464514 265618 464546 265854
rect 464782 265618 464866 265854
rect 465102 265618 465134 265854
rect 464514 226174 465134 265618
rect 464514 225938 464546 226174
rect 464782 225938 464866 226174
rect 465102 225938 465134 226174
rect 464514 225854 465134 225938
rect 464514 225618 464546 225854
rect 464782 225618 464866 225854
rect 465102 225618 465134 225854
rect 464514 186174 465134 225618
rect 464514 185938 464546 186174
rect 464782 185938 464866 186174
rect 465102 185938 465134 186174
rect 464514 185854 465134 185938
rect 464514 185618 464546 185854
rect 464782 185618 464866 185854
rect 465102 185618 465134 185854
rect 464514 146174 465134 185618
rect 464514 145938 464546 146174
rect 464782 145938 464866 146174
rect 465102 145938 465134 146174
rect 464514 145854 465134 145938
rect 464514 145618 464546 145854
rect 464782 145618 464866 145854
rect 465102 145618 465134 145854
rect 464514 106174 465134 145618
rect 464514 105938 464546 106174
rect 464782 105938 464866 106174
rect 465102 105938 465134 106174
rect 464514 105854 465134 105938
rect 464514 105618 464546 105854
rect 464782 105618 464866 105854
rect 465102 105618 465134 105854
rect 464514 66174 465134 105618
rect 464514 65938 464546 66174
rect 464782 65938 464866 66174
rect 465102 65938 465134 66174
rect 464514 65854 465134 65938
rect 464514 65618 464546 65854
rect 464782 65618 464866 65854
rect 465102 65618 465134 65854
rect 464514 26174 465134 65618
rect 464514 25938 464546 26174
rect 464782 25938 464866 26174
rect 465102 25938 465134 26174
rect 464514 25854 465134 25938
rect 464514 25618 464546 25854
rect 464782 25618 464866 25854
rect 465102 25618 465134 25854
rect 464514 -3226 465134 25618
rect 464514 -3462 464546 -3226
rect 464782 -3462 464866 -3226
rect 465102 -3462 465134 -3226
rect 464514 -3546 465134 -3462
rect 464514 -3782 464546 -3546
rect 464782 -3782 464866 -3546
rect 465102 -3782 465134 -3546
rect 464514 -3814 465134 -3782
rect 468234 669894 468854 709082
rect 468234 669658 468266 669894
rect 468502 669658 468586 669894
rect 468822 669658 468854 669894
rect 468234 669574 468854 669658
rect 468234 669338 468266 669574
rect 468502 669338 468586 669574
rect 468822 669338 468854 669574
rect 468234 629894 468854 669338
rect 468234 629658 468266 629894
rect 468502 629658 468586 629894
rect 468822 629658 468854 629894
rect 468234 629574 468854 629658
rect 468234 629338 468266 629574
rect 468502 629338 468586 629574
rect 468822 629338 468854 629574
rect 468234 589894 468854 629338
rect 468234 589658 468266 589894
rect 468502 589658 468586 589894
rect 468822 589658 468854 589894
rect 468234 589574 468854 589658
rect 468234 589338 468266 589574
rect 468502 589338 468586 589574
rect 468822 589338 468854 589574
rect 468234 549894 468854 589338
rect 468234 549658 468266 549894
rect 468502 549658 468586 549894
rect 468822 549658 468854 549894
rect 468234 549574 468854 549658
rect 468234 549338 468266 549574
rect 468502 549338 468586 549574
rect 468822 549338 468854 549574
rect 468234 509894 468854 549338
rect 468234 509658 468266 509894
rect 468502 509658 468586 509894
rect 468822 509658 468854 509894
rect 468234 509574 468854 509658
rect 468234 509338 468266 509574
rect 468502 509338 468586 509574
rect 468822 509338 468854 509574
rect 468234 469894 468854 509338
rect 468234 469658 468266 469894
rect 468502 469658 468586 469894
rect 468822 469658 468854 469894
rect 468234 469574 468854 469658
rect 468234 469338 468266 469574
rect 468502 469338 468586 469574
rect 468822 469338 468854 469574
rect 468234 429894 468854 469338
rect 468234 429658 468266 429894
rect 468502 429658 468586 429894
rect 468822 429658 468854 429894
rect 468234 429574 468854 429658
rect 468234 429338 468266 429574
rect 468502 429338 468586 429574
rect 468822 429338 468854 429574
rect 468234 389894 468854 429338
rect 468234 389658 468266 389894
rect 468502 389658 468586 389894
rect 468822 389658 468854 389894
rect 468234 389574 468854 389658
rect 468234 389338 468266 389574
rect 468502 389338 468586 389574
rect 468822 389338 468854 389574
rect 468234 349894 468854 389338
rect 468234 349658 468266 349894
rect 468502 349658 468586 349894
rect 468822 349658 468854 349894
rect 468234 349574 468854 349658
rect 468234 349338 468266 349574
rect 468502 349338 468586 349574
rect 468822 349338 468854 349574
rect 468234 309894 468854 349338
rect 468234 309658 468266 309894
rect 468502 309658 468586 309894
rect 468822 309658 468854 309894
rect 468234 309574 468854 309658
rect 468234 309338 468266 309574
rect 468502 309338 468586 309574
rect 468822 309338 468854 309574
rect 468234 269894 468854 309338
rect 468234 269658 468266 269894
rect 468502 269658 468586 269894
rect 468822 269658 468854 269894
rect 468234 269574 468854 269658
rect 468234 269338 468266 269574
rect 468502 269338 468586 269574
rect 468822 269338 468854 269574
rect 468234 229894 468854 269338
rect 468234 229658 468266 229894
rect 468502 229658 468586 229894
rect 468822 229658 468854 229894
rect 468234 229574 468854 229658
rect 468234 229338 468266 229574
rect 468502 229338 468586 229574
rect 468822 229338 468854 229574
rect 468234 189894 468854 229338
rect 468234 189658 468266 189894
rect 468502 189658 468586 189894
rect 468822 189658 468854 189894
rect 468234 189574 468854 189658
rect 468234 189338 468266 189574
rect 468502 189338 468586 189574
rect 468822 189338 468854 189574
rect 468234 149894 468854 189338
rect 468234 149658 468266 149894
rect 468502 149658 468586 149894
rect 468822 149658 468854 149894
rect 468234 149574 468854 149658
rect 468234 149338 468266 149574
rect 468502 149338 468586 149574
rect 468822 149338 468854 149574
rect 468234 109894 468854 149338
rect 468234 109658 468266 109894
rect 468502 109658 468586 109894
rect 468822 109658 468854 109894
rect 468234 109574 468854 109658
rect 468234 109338 468266 109574
rect 468502 109338 468586 109574
rect 468822 109338 468854 109574
rect 468234 69894 468854 109338
rect 468234 69658 468266 69894
rect 468502 69658 468586 69894
rect 468822 69658 468854 69894
rect 468234 69574 468854 69658
rect 468234 69338 468266 69574
rect 468502 69338 468586 69574
rect 468822 69338 468854 69574
rect 468234 29894 468854 69338
rect 468234 29658 468266 29894
rect 468502 29658 468586 29894
rect 468822 29658 468854 29894
rect 468234 29574 468854 29658
rect 468234 29338 468266 29574
rect 468502 29338 468586 29574
rect 468822 29338 468854 29574
rect 468234 -5146 468854 29338
rect 468234 -5382 468266 -5146
rect 468502 -5382 468586 -5146
rect 468822 -5382 468854 -5146
rect 468234 -5466 468854 -5382
rect 468234 -5702 468266 -5466
rect 468502 -5702 468586 -5466
rect 468822 -5702 468854 -5466
rect 468234 -5734 468854 -5702
rect 471954 673614 472574 711002
rect 491954 710598 492574 711590
rect 491954 710362 491986 710598
rect 492222 710362 492306 710598
rect 492542 710362 492574 710598
rect 491954 710278 492574 710362
rect 491954 710042 491986 710278
rect 492222 710042 492306 710278
rect 492542 710042 492574 710278
rect 488234 708678 488854 709670
rect 488234 708442 488266 708678
rect 488502 708442 488586 708678
rect 488822 708442 488854 708678
rect 488234 708358 488854 708442
rect 488234 708122 488266 708358
rect 488502 708122 488586 708358
rect 488822 708122 488854 708358
rect 484514 706758 485134 707750
rect 484514 706522 484546 706758
rect 484782 706522 484866 706758
rect 485102 706522 485134 706758
rect 484514 706438 485134 706522
rect 484514 706202 484546 706438
rect 484782 706202 484866 706438
rect 485102 706202 485134 706438
rect 471954 673378 471986 673614
rect 472222 673378 472306 673614
rect 472542 673378 472574 673614
rect 471954 673294 472574 673378
rect 471954 673058 471986 673294
rect 472222 673058 472306 673294
rect 472542 673058 472574 673294
rect 471954 633614 472574 673058
rect 471954 633378 471986 633614
rect 472222 633378 472306 633614
rect 472542 633378 472574 633614
rect 471954 633294 472574 633378
rect 471954 633058 471986 633294
rect 472222 633058 472306 633294
rect 472542 633058 472574 633294
rect 471954 593614 472574 633058
rect 471954 593378 471986 593614
rect 472222 593378 472306 593614
rect 472542 593378 472574 593614
rect 471954 593294 472574 593378
rect 471954 593058 471986 593294
rect 472222 593058 472306 593294
rect 472542 593058 472574 593294
rect 471954 553614 472574 593058
rect 471954 553378 471986 553614
rect 472222 553378 472306 553614
rect 472542 553378 472574 553614
rect 471954 553294 472574 553378
rect 471954 553058 471986 553294
rect 472222 553058 472306 553294
rect 472542 553058 472574 553294
rect 471954 513614 472574 553058
rect 471954 513378 471986 513614
rect 472222 513378 472306 513614
rect 472542 513378 472574 513614
rect 471954 513294 472574 513378
rect 471954 513058 471986 513294
rect 472222 513058 472306 513294
rect 472542 513058 472574 513294
rect 471954 473614 472574 513058
rect 471954 473378 471986 473614
rect 472222 473378 472306 473614
rect 472542 473378 472574 473614
rect 471954 473294 472574 473378
rect 471954 473058 471986 473294
rect 472222 473058 472306 473294
rect 472542 473058 472574 473294
rect 471954 433614 472574 473058
rect 471954 433378 471986 433614
rect 472222 433378 472306 433614
rect 472542 433378 472574 433614
rect 471954 433294 472574 433378
rect 471954 433058 471986 433294
rect 472222 433058 472306 433294
rect 472542 433058 472574 433294
rect 471954 393614 472574 433058
rect 471954 393378 471986 393614
rect 472222 393378 472306 393614
rect 472542 393378 472574 393614
rect 471954 393294 472574 393378
rect 471954 393058 471986 393294
rect 472222 393058 472306 393294
rect 472542 393058 472574 393294
rect 471954 353614 472574 393058
rect 471954 353378 471986 353614
rect 472222 353378 472306 353614
rect 472542 353378 472574 353614
rect 471954 353294 472574 353378
rect 471954 353058 471986 353294
rect 472222 353058 472306 353294
rect 472542 353058 472574 353294
rect 471954 313614 472574 353058
rect 471954 313378 471986 313614
rect 472222 313378 472306 313614
rect 472542 313378 472574 313614
rect 471954 313294 472574 313378
rect 471954 313058 471986 313294
rect 472222 313058 472306 313294
rect 472542 313058 472574 313294
rect 471954 273614 472574 313058
rect 471954 273378 471986 273614
rect 472222 273378 472306 273614
rect 472542 273378 472574 273614
rect 471954 273294 472574 273378
rect 471954 273058 471986 273294
rect 472222 273058 472306 273294
rect 472542 273058 472574 273294
rect 471954 233614 472574 273058
rect 471954 233378 471986 233614
rect 472222 233378 472306 233614
rect 472542 233378 472574 233614
rect 471954 233294 472574 233378
rect 471954 233058 471986 233294
rect 472222 233058 472306 233294
rect 472542 233058 472574 233294
rect 471954 193614 472574 233058
rect 471954 193378 471986 193614
rect 472222 193378 472306 193614
rect 472542 193378 472574 193614
rect 471954 193294 472574 193378
rect 471954 193058 471986 193294
rect 472222 193058 472306 193294
rect 472542 193058 472574 193294
rect 471954 153614 472574 193058
rect 471954 153378 471986 153614
rect 472222 153378 472306 153614
rect 472542 153378 472574 153614
rect 471954 153294 472574 153378
rect 471954 153058 471986 153294
rect 472222 153058 472306 153294
rect 472542 153058 472574 153294
rect 471954 113614 472574 153058
rect 471954 113378 471986 113614
rect 472222 113378 472306 113614
rect 472542 113378 472574 113614
rect 471954 113294 472574 113378
rect 471954 113058 471986 113294
rect 472222 113058 472306 113294
rect 472542 113058 472574 113294
rect 471954 73614 472574 113058
rect 471954 73378 471986 73614
rect 472222 73378 472306 73614
rect 472542 73378 472574 73614
rect 471954 73294 472574 73378
rect 471954 73058 471986 73294
rect 472222 73058 472306 73294
rect 472542 73058 472574 73294
rect 471954 33614 472574 73058
rect 471954 33378 471986 33614
rect 472222 33378 472306 33614
rect 472542 33378 472574 33614
rect 471954 33294 472574 33378
rect 471954 33058 471986 33294
rect 472222 33058 472306 33294
rect 472542 33058 472574 33294
rect 451954 -6342 451986 -6106
rect 452222 -6342 452306 -6106
rect 452542 -6342 452574 -6106
rect 451954 -6426 452574 -6342
rect 451954 -6662 451986 -6426
rect 452222 -6662 452306 -6426
rect 452542 -6662 452574 -6426
rect 451954 -7654 452574 -6662
rect 471954 -7066 472574 33058
rect 480794 704838 481414 705830
rect 480794 704602 480826 704838
rect 481062 704602 481146 704838
rect 481382 704602 481414 704838
rect 480794 704518 481414 704602
rect 480794 704282 480826 704518
rect 481062 704282 481146 704518
rect 481382 704282 481414 704518
rect 480794 682454 481414 704282
rect 480794 682218 480826 682454
rect 481062 682218 481146 682454
rect 481382 682218 481414 682454
rect 480794 682134 481414 682218
rect 480794 681898 480826 682134
rect 481062 681898 481146 682134
rect 481382 681898 481414 682134
rect 480794 642454 481414 681898
rect 480794 642218 480826 642454
rect 481062 642218 481146 642454
rect 481382 642218 481414 642454
rect 480794 642134 481414 642218
rect 480794 641898 480826 642134
rect 481062 641898 481146 642134
rect 481382 641898 481414 642134
rect 480794 602454 481414 641898
rect 480794 602218 480826 602454
rect 481062 602218 481146 602454
rect 481382 602218 481414 602454
rect 480794 602134 481414 602218
rect 480794 601898 480826 602134
rect 481062 601898 481146 602134
rect 481382 601898 481414 602134
rect 480794 562454 481414 601898
rect 480794 562218 480826 562454
rect 481062 562218 481146 562454
rect 481382 562218 481414 562454
rect 480794 562134 481414 562218
rect 480794 561898 480826 562134
rect 481062 561898 481146 562134
rect 481382 561898 481414 562134
rect 480794 522454 481414 561898
rect 480794 522218 480826 522454
rect 481062 522218 481146 522454
rect 481382 522218 481414 522454
rect 480794 522134 481414 522218
rect 480794 521898 480826 522134
rect 481062 521898 481146 522134
rect 481382 521898 481414 522134
rect 480794 482454 481414 521898
rect 480794 482218 480826 482454
rect 481062 482218 481146 482454
rect 481382 482218 481414 482454
rect 480794 482134 481414 482218
rect 480794 481898 480826 482134
rect 481062 481898 481146 482134
rect 481382 481898 481414 482134
rect 480794 442454 481414 481898
rect 480794 442218 480826 442454
rect 481062 442218 481146 442454
rect 481382 442218 481414 442454
rect 480794 442134 481414 442218
rect 480794 441898 480826 442134
rect 481062 441898 481146 442134
rect 481382 441898 481414 442134
rect 480794 402454 481414 441898
rect 480794 402218 480826 402454
rect 481062 402218 481146 402454
rect 481382 402218 481414 402454
rect 480794 402134 481414 402218
rect 480794 401898 480826 402134
rect 481062 401898 481146 402134
rect 481382 401898 481414 402134
rect 480794 362454 481414 401898
rect 480794 362218 480826 362454
rect 481062 362218 481146 362454
rect 481382 362218 481414 362454
rect 480794 362134 481414 362218
rect 480794 361898 480826 362134
rect 481062 361898 481146 362134
rect 481382 361898 481414 362134
rect 480794 322454 481414 361898
rect 480794 322218 480826 322454
rect 481062 322218 481146 322454
rect 481382 322218 481414 322454
rect 480794 322134 481414 322218
rect 480794 321898 480826 322134
rect 481062 321898 481146 322134
rect 481382 321898 481414 322134
rect 480794 282454 481414 321898
rect 480794 282218 480826 282454
rect 481062 282218 481146 282454
rect 481382 282218 481414 282454
rect 480794 282134 481414 282218
rect 480794 281898 480826 282134
rect 481062 281898 481146 282134
rect 481382 281898 481414 282134
rect 480794 242454 481414 281898
rect 480794 242218 480826 242454
rect 481062 242218 481146 242454
rect 481382 242218 481414 242454
rect 480794 242134 481414 242218
rect 480794 241898 480826 242134
rect 481062 241898 481146 242134
rect 481382 241898 481414 242134
rect 480794 202454 481414 241898
rect 480794 202218 480826 202454
rect 481062 202218 481146 202454
rect 481382 202218 481414 202454
rect 480794 202134 481414 202218
rect 480794 201898 480826 202134
rect 481062 201898 481146 202134
rect 481382 201898 481414 202134
rect 480794 162454 481414 201898
rect 480794 162218 480826 162454
rect 481062 162218 481146 162454
rect 481382 162218 481414 162454
rect 480794 162134 481414 162218
rect 480794 161898 480826 162134
rect 481062 161898 481146 162134
rect 481382 161898 481414 162134
rect 480794 122454 481414 161898
rect 480794 122218 480826 122454
rect 481062 122218 481146 122454
rect 481382 122218 481414 122454
rect 480794 122134 481414 122218
rect 480794 121898 480826 122134
rect 481062 121898 481146 122134
rect 481382 121898 481414 122134
rect 480794 82454 481414 121898
rect 480794 82218 480826 82454
rect 481062 82218 481146 82454
rect 481382 82218 481414 82454
rect 480794 82134 481414 82218
rect 480794 81898 480826 82134
rect 481062 81898 481146 82134
rect 481382 81898 481414 82134
rect 480794 42454 481414 81898
rect 480794 42218 480826 42454
rect 481062 42218 481146 42454
rect 481382 42218 481414 42454
rect 480794 42134 481414 42218
rect 480794 41898 480826 42134
rect 481062 41898 481146 42134
rect 481382 41898 481414 42134
rect 480794 2454 481414 41898
rect 480794 2218 480826 2454
rect 481062 2218 481146 2454
rect 481382 2218 481414 2454
rect 480794 2134 481414 2218
rect 480794 1898 480826 2134
rect 481062 1898 481146 2134
rect 481382 1898 481414 2134
rect 480794 -346 481414 1898
rect 480794 -582 480826 -346
rect 481062 -582 481146 -346
rect 481382 -582 481414 -346
rect 480794 -666 481414 -582
rect 480794 -902 480826 -666
rect 481062 -902 481146 -666
rect 481382 -902 481414 -666
rect 480794 -1894 481414 -902
rect 484514 686174 485134 706202
rect 484514 685938 484546 686174
rect 484782 685938 484866 686174
rect 485102 685938 485134 686174
rect 484514 685854 485134 685938
rect 484514 685618 484546 685854
rect 484782 685618 484866 685854
rect 485102 685618 485134 685854
rect 484514 646174 485134 685618
rect 484514 645938 484546 646174
rect 484782 645938 484866 646174
rect 485102 645938 485134 646174
rect 484514 645854 485134 645938
rect 484514 645618 484546 645854
rect 484782 645618 484866 645854
rect 485102 645618 485134 645854
rect 484514 606174 485134 645618
rect 484514 605938 484546 606174
rect 484782 605938 484866 606174
rect 485102 605938 485134 606174
rect 484514 605854 485134 605938
rect 484514 605618 484546 605854
rect 484782 605618 484866 605854
rect 485102 605618 485134 605854
rect 484514 566174 485134 605618
rect 484514 565938 484546 566174
rect 484782 565938 484866 566174
rect 485102 565938 485134 566174
rect 484514 565854 485134 565938
rect 484514 565618 484546 565854
rect 484782 565618 484866 565854
rect 485102 565618 485134 565854
rect 484514 526174 485134 565618
rect 484514 525938 484546 526174
rect 484782 525938 484866 526174
rect 485102 525938 485134 526174
rect 484514 525854 485134 525938
rect 484514 525618 484546 525854
rect 484782 525618 484866 525854
rect 485102 525618 485134 525854
rect 484514 486174 485134 525618
rect 484514 485938 484546 486174
rect 484782 485938 484866 486174
rect 485102 485938 485134 486174
rect 484514 485854 485134 485938
rect 484514 485618 484546 485854
rect 484782 485618 484866 485854
rect 485102 485618 485134 485854
rect 484514 446174 485134 485618
rect 484514 445938 484546 446174
rect 484782 445938 484866 446174
rect 485102 445938 485134 446174
rect 484514 445854 485134 445938
rect 484514 445618 484546 445854
rect 484782 445618 484866 445854
rect 485102 445618 485134 445854
rect 484514 406174 485134 445618
rect 484514 405938 484546 406174
rect 484782 405938 484866 406174
rect 485102 405938 485134 406174
rect 484514 405854 485134 405938
rect 484514 405618 484546 405854
rect 484782 405618 484866 405854
rect 485102 405618 485134 405854
rect 484514 366174 485134 405618
rect 484514 365938 484546 366174
rect 484782 365938 484866 366174
rect 485102 365938 485134 366174
rect 484514 365854 485134 365938
rect 484514 365618 484546 365854
rect 484782 365618 484866 365854
rect 485102 365618 485134 365854
rect 484514 326174 485134 365618
rect 484514 325938 484546 326174
rect 484782 325938 484866 326174
rect 485102 325938 485134 326174
rect 484514 325854 485134 325938
rect 484514 325618 484546 325854
rect 484782 325618 484866 325854
rect 485102 325618 485134 325854
rect 484514 286174 485134 325618
rect 484514 285938 484546 286174
rect 484782 285938 484866 286174
rect 485102 285938 485134 286174
rect 484514 285854 485134 285938
rect 484514 285618 484546 285854
rect 484782 285618 484866 285854
rect 485102 285618 485134 285854
rect 484514 246174 485134 285618
rect 484514 245938 484546 246174
rect 484782 245938 484866 246174
rect 485102 245938 485134 246174
rect 484514 245854 485134 245938
rect 484514 245618 484546 245854
rect 484782 245618 484866 245854
rect 485102 245618 485134 245854
rect 484514 206174 485134 245618
rect 484514 205938 484546 206174
rect 484782 205938 484866 206174
rect 485102 205938 485134 206174
rect 484514 205854 485134 205938
rect 484514 205618 484546 205854
rect 484782 205618 484866 205854
rect 485102 205618 485134 205854
rect 484514 166174 485134 205618
rect 484514 165938 484546 166174
rect 484782 165938 484866 166174
rect 485102 165938 485134 166174
rect 484514 165854 485134 165938
rect 484514 165618 484546 165854
rect 484782 165618 484866 165854
rect 485102 165618 485134 165854
rect 484514 126174 485134 165618
rect 484514 125938 484546 126174
rect 484782 125938 484866 126174
rect 485102 125938 485134 126174
rect 484514 125854 485134 125938
rect 484514 125618 484546 125854
rect 484782 125618 484866 125854
rect 485102 125618 485134 125854
rect 484514 86174 485134 125618
rect 484514 85938 484546 86174
rect 484782 85938 484866 86174
rect 485102 85938 485134 86174
rect 484514 85854 485134 85938
rect 484514 85618 484546 85854
rect 484782 85618 484866 85854
rect 485102 85618 485134 85854
rect 484514 46174 485134 85618
rect 484514 45938 484546 46174
rect 484782 45938 484866 46174
rect 485102 45938 485134 46174
rect 484514 45854 485134 45938
rect 484514 45618 484546 45854
rect 484782 45618 484866 45854
rect 485102 45618 485134 45854
rect 484514 6174 485134 45618
rect 484514 5938 484546 6174
rect 484782 5938 484866 6174
rect 485102 5938 485134 6174
rect 484514 5854 485134 5938
rect 484514 5618 484546 5854
rect 484782 5618 484866 5854
rect 485102 5618 485134 5854
rect 484514 -2266 485134 5618
rect 484514 -2502 484546 -2266
rect 484782 -2502 484866 -2266
rect 485102 -2502 485134 -2266
rect 484514 -2586 485134 -2502
rect 484514 -2822 484546 -2586
rect 484782 -2822 484866 -2586
rect 485102 -2822 485134 -2586
rect 484514 -3814 485134 -2822
rect 488234 689894 488854 708122
rect 488234 689658 488266 689894
rect 488502 689658 488586 689894
rect 488822 689658 488854 689894
rect 488234 689574 488854 689658
rect 488234 689338 488266 689574
rect 488502 689338 488586 689574
rect 488822 689338 488854 689574
rect 488234 649894 488854 689338
rect 488234 649658 488266 649894
rect 488502 649658 488586 649894
rect 488822 649658 488854 649894
rect 488234 649574 488854 649658
rect 488234 649338 488266 649574
rect 488502 649338 488586 649574
rect 488822 649338 488854 649574
rect 488234 609894 488854 649338
rect 488234 609658 488266 609894
rect 488502 609658 488586 609894
rect 488822 609658 488854 609894
rect 488234 609574 488854 609658
rect 488234 609338 488266 609574
rect 488502 609338 488586 609574
rect 488822 609338 488854 609574
rect 488234 569894 488854 609338
rect 488234 569658 488266 569894
rect 488502 569658 488586 569894
rect 488822 569658 488854 569894
rect 488234 569574 488854 569658
rect 488234 569338 488266 569574
rect 488502 569338 488586 569574
rect 488822 569338 488854 569574
rect 488234 529894 488854 569338
rect 488234 529658 488266 529894
rect 488502 529658 488586 529894
rect 488822 529658 488854 529894
rect 488234 529574 488854 529658
rect 488234 529338 488266 529574
rect 488502 529338 488586 529574
rect 488822 529338 488854 529574
rect 488234 489894 488854 529338
rect 488234 489658 488266 489894
rect 488502 489658 488586 489894
rect 488822 489658 488854 489894
rect 488234 489574 488854 489658
rect 488234 489338 488266 489574
rect 488502 489338 488586 489574
rect 488822 489338 488854 489574
rect 488234 449894 488854 489338
rect 488234 449658 488266 449894
rect 488502 449658 488586 449894
rect 488822 449658 488854 449894
rect 488234 449574 488854 449658
rect 488234 449338 488266 449574
rect 488502 449338 488586 449574
rect 488822 449338 488854 449574
rect 488234 409894 488854 449338
rect 488234 409658 488266 409894
rect 488502 409658 488586 409894
rect 488822 409658 488854 409894
rect 488234 409574 488854 409658
rect 488234 409338 488266 409574
rect 488502 409338 488586 409574
rect 488822 409338 488854 409574
rect 488234 369894 488854 409338
rect 488234 369658 488266 369894
rect 488502 369658 488586 369894
rect 488822 369658 488854 369894
rect 488234 369574 488854 369658
rect 488234 369338 488266 369574
rect 488502 369338 488586 369574
rect 488822 369338 488854 369574
rect 488234 329894 488854 369338
rect 488234 329658 488266 329894
rect 488502 329658 488586 329894
rect 488822 329658 488854 329894
rect 488234 329574 488854 329658
rect 488234 329338 488266 329574
rect 488502 329338 488586 329574
rect 488822 329338 488854 329574
rect 488234 289894 488854 329338
rect 488234 289658 488266 289894
rect 488502 289658 488586 289894
rect 488822 289658 488854 289894
rect 488234 289574 488854 289658
rect 488234 289338 488266 289574
rect 488502 289338 488586 289574
rect 488822 289338 488854 289574
rect 488234 249894 488854 289338
rect 488234 249658 488266 249894
rect 488502 249658 488586 249894
rect 488822 249658 488854 249894
rect 488234 249574 488854 249658
rect 488234 249338 488266 249574
rect 488502 249338 488586 249574
rect 488822 249338 488854 249574
rect 488234 209894 488854 249338
rect 488234 209658 488266 209894
rect 488502 209658 488586 209894
rect 488822 209658 488854 209894
rect 488234 209574 488854 209658
rect 488234 209338 488266 209574
rect 488502 209338 488586 209574
rect 488822 209338 488854 209574
rect 488234 169894 488854 209338
rect 488234 169658 488266 169894
rect 488502 169658 488586 169894
rect 488822 169658 488854 169894
rect 488234 169574 488854 169658
rect 488234 169338 488266 169574
rect 488502 169338 488586 169574
rect 488822 169338 488854 169574
rect 488234 129894 488854 169338
rect 488234 129658 488266 129894
rect 488502 129658 488586 129894
rect 488822 129658 488854 129894
rect 488234 129574 488854 129658
rect 488234 129338 488266 129574
rect 488502 129338 488586 129574
rect 488822 129338 488854 129574
rect 488234 89894 488854 129338
rect 488234 89658 488266 89894
rect 488502 89658 488586 89894
rect 488822 89658 488854 89894
rect 488234 89574 488854 89658
rect 488234 89338 488266 89574
rect 488502 89338 488586 89574
rect 488822 89338 488854 89574
rect 488234 49894 488854 89338
rect 488234 49658 488266 49894
rect 488502 49658 488586 49894
rect 488822 49658 488854 49894
rect 488234 49574 488854 49658
rect 488234 49338 488266 49574
rect 488502 49338 488586 49574
rect 488822 49338 488854 49574
rect 488234 9894 488854 49338
rect 488234 9658 488266 9894
rect 488502 9658 488586 9894
rect 488822 9658 488854 9894
rect 488234 9574 488854 9658
rect 488234 9338 488266 9574
rect 488502 9338 488586 9574
rect 488822 9338 488854 9574
rect 488234 -4186 488854 9338
rect 488234 -4422 488266 -4186
rect 488502 -4422 488586 -4186
rect 488822 -4422 488854 -4186
rect 488234 -4506 488854 -4422
rect 488234 -4742 488266 -4506
rect 488502 -4742 488586 -4506
rect 488822 -4742 488854 -4506
rect 488234 -5734 488854 -4742
rect 491954 693614 492574 710042
rect 511954 711558 512574 711590
rect 511954 711322 511986 711558
rect 512222 711322 512306 711558
rect 512542 711322 512574 711558
rect 511954 711238 512574 711322
rect 511954 711002 511986 711238
rect 512222 711002 512306 711238
rect 512542 711002 512574 711238
rect 508234 709638 508854 709670
rect 508234 709402 508266 709638
rect 508502 709402 508586 709638
rect 508822 709402 508854 709638
rect 508234 709318 508854 709402
rect 508234 709082 508266 709318
rect 508502 709082 508586 709318
rect 508822 709082 508854 709318
rect 504514 707718 505134 707750
rect 504514 707482 504546 707718
rect 504782 707482 504866 707718
rect 505102 707482 505134 707718
rect 504514 707398 505134 707482
rect 504514 707162 504546 707398
rect 504782 707162 504866 707398
rect 505102 707162 505134 707398
rect 491954 693378 491986 693614
rect 492222 693378 492306 693614
rect 492542 693378 492574 693614
rect 491954 693294 492574 693378
rect 491954 693058 491986 693294
rect 492222 693058 492306 693294
rect 492542 693058 492574 693294
rect 491954 653614 492574 693058
rect 491954 653378 491986 653614
rect 492222 653378 492306 653614
rect 492542 653378 492574 653614
rect 491954 653294 492574 653378
rect 491954 653058 491986 653294
rect 492222 653058 492306 653294
rect 492542 653058 492574 653294
rect 491954 613614 492574 653058
rect 491954 613378 491986 613614
rect 492222 613378 492306 613614
rect 492542 613378 492574 613614
rect 491954 613294 492574 613378
rect 491954 613058 491986 613294
rect 492222 613058 492306 613294
rect 492542 613058 492574 613294
rect 491954 573614 492574 613058
rect 491954 573378 491986 573614
rect 492222 573378 492306 573614
rect 492542 573378 492574 573614
rect 491954 573294 492574 573378
rect 491954 573058 491986 573294
rect 492222 573058 492306 573294
rect 492542 573058 492574 573294
rect 491954 533614 492574 573058
rect 491954 533378 491986 533614
rect 492222 533378 492306 533614
rect 492542 533378 492574 533614
rect 491954 533294 492574 533378
rect 491954 533058 491986 533294
rect 492222 533058 492306 533294
rect 492542 533058 492574 533294
rect 491954 493614 492574 533058
rect 491954 493378 491986 493614
rect 492222 493378 492306 493614
rect 492542 493378 492574 493614
rect 491954 493294 492574 493378
rect 491954 493058 491986 493294
rect 492222 493058 492306 493294
rect 492542 493058 492574 493294
rect 491954 453614 492574 493058
rect 491954 453378 491986 453614
rect 492222 453378 492306 453614
rect 492542 453378 492574 453614
rect 491954 453294 492574 453378
rect 491954 453058 491986 453294
rect 492222 453058 492306 453294
rect 492542 453058 492574 453294
rect 491954 413614 492574 453058
rect 491954 413378 491986 413614
rect 492222 413378 492306 413614
rect 492542 413378 492574 413614
rect 491954 413294 492574 413378
rect 491954 413058 491986 413294
rect 492222 413058 492306 413294
rect 492542 413058 492574 413294
rect 491954 373614 492574 413058
rect 491954 373378 491986 373614
rect 492222 373378 492306 373614
rect 492542 373378 492574 373614
rect 491954 373294 492574 373378
rect 491954 373058 491986 373294
rect 492222 373058 492306 373294
rect 492542 373058 492574 373294
rect 491954 333614 492574 373058
rect 491954 333378 491986 333614
rect 492222 333378 492306 333614
rect 492542 333378 492574 333614
rect 491954 333294 492574 333378
rect 491954 333058 491986 333294
rect 492222 333058 492306 333294
rect 492542 333058 492574 333294
rect 491954 293614 492574 333058
rect 491954 293378 491986 293614
rect 492222 293378 492306 293614
rect 492542 293378 492574 293614
rect 491954 293294 492574 293378
rect 491954 293058 491986 293294
rect 492222 293058 492306 293294
rect 492542 293058 492574 293294
rect 491954 253614 492574 293058
rect 491954 253378 491986 253614
rect 492222 253378 492306 253614
rect 492542 253378 492574 253614
rect 491954 253294 492574 253378
rect 491954 253058 491986 253294
rect 492222 253058 492306 253294
rect 492542 253058 492574 253294
rect 491954 213614 492574 253058
rect 491954 213378 491986 213614
rect 492222 213378 492306 213614
rect 492542 213378 492574 213614
rect 491954 213294 492574 213378
rect 491954 213058 491986 213294
rect 492222 213058 492306 213294
rect 492542 213058 492574 213294
rect 491954 173614 492574 213058
rect 491954 173378 491986 173614
rect 492222 173378 492306 173614
rect 492542 173378 492574 173614
rect 491954 173294 492574 173378
rect 491954 173058 491986 173294
rect 492222 173058 492306 173294
rect 492542 173058 492574 173294
rect 491954 133614 492574 173058
rect 491954 133378 491986 133614
rect 492222 133378 492306 133614
rect 492542 133378 492574 133614
rect 491954 133294 492574 133378
rect 491954 133058 491986 133294
rect 492222 133058 492306 133294
rect 492542 133058 492574 133294
rect 491954 93614 492574 133058
rect 491954 93378 491986 93614
rect 492222 93378 492306 93614
rect 492542 93378 492574 93614
rect 491954 93294 492574 93378
rect 491954 93058 491986 93294
rect 492222 93058 492306 93294
rect 492542 93058 492574 93294
rect 491954 53614 492574 93058
rect 491954 53378 491986 53614
rect 492222 53378 492306 53614
rect 492542 53378 492574 53614
rect 491954 53294 492574 53378
rect 491954 53058 491986 53294
rect 492222 53058 492306 53294
rect 492542 53058 492574 53294
rect 491954 13614 492574 53058
rect 491954 13378 491986 13614
rect 492222 13378 492306 13614
rect 492542 13378 492574 13614
rect 491954 13294 492574 13378
rect 491954 13058 491986 13294
rect 492222 13058 492306 13294
rect 492542 13058 492574 13294
rect 471954 -7302 471986 -7066
rect 472222 -7302 472306 -7066
rect 472542 -7302 472574 -7066
rect 471954 -7386 472574 -7302
rect 471954 -7622 471986 -7386
rect 472222 -7622 472306 -7386
rect 472542 -7622 472574 -7386
rect 471954 -7654 472574 -7622
rect 491954 -6106 492574 13058
rect 500794 705798 501414 705830
rect 500794 705562 500826 705798
rect 501062 705562 501146 705798
rect 501382 705562 501414 705798
rect 500794 705478 501414 705562
rect 500794 705242 500826 705478
rect 501062 705242 501146 705478
rect 501382 705242 501414 705478
rect 500794 662454 501414 705242
rect 500794 662218 500826 662454
rect 501062 662218 501146 662454
rect 501382 662218 501414 662454
rect 500794 662134 501414 662218
rect 500794 661898 500826 662134
rect 501062 661898 501146 662134
rect 501382 661898 501414 662134
rect 500794 622454 501414 661898
rect 500794 622218 500826 622454
rect 501062 622218 501146 622454
rect 501382 622218 501414 622454
rect 500794 622134 501414 622218
rect 500794 621898 500826 622134
rect 501062 621898 501146 622134
rect 501382 621898 501414 622134
rect 500794 582454 501414 621898
rect 500794 582218 500826 582454
rect 501062 582218 501146 582454
rect 501382 582218 501414 582454
rect 500794 582134 501414 582218
rect 500794 581898 500826 582134
rect 501062 581898 501146 582134
rect 501382 581898 501414 582134
rect 500794 542454 501414 581898
rect 500794 542218 500826 542454
rect 501062 542218 501146 542454
rect 501382 542218 501414 542454
rect 500794 542134 501414 542218
rect 500794 541898 500826 542134
rect 501062 541898 501146 542134
rect 501382 541898 501414 542134
rect 500794 502454 501414 541898
rect 500794 502218 500826 502454
rect 501062 502218 501146 502454
rect 501382 502218 501414 502454
rect 500794 502134 501414 502218
rect 500794 501898 500826 502134
rect 501062 501898 501146 502134
rect 501382 501898 501414 502134
rect 500794 462454 501414 501898
rect 500794 462218 500826 462454
rect 501062 462218 501146 462454
rect 501382 462218 501414 462454
rect 500794 462134 501414 462218
rect 500794 461898 500826 462134
rect 501062 461898 501146 462134
rect 501382 461898 501414 462134
rect 500794 422454 501414 461898
rect 500794 422218 500826 422454
rect 501062 422218 501146 422454
rect 501382 422218 501414 422454
rect 500794 422134 501414 422218
rect 500794 421898 500826 422134
rect 501062 421898 501146 422134
rect 501382 421898 501414 422134
rect 500794 382454 501414 421898
rect 500794 382218 500826 382454
rect 501062 382218 501146 382454
rect 501382 382218 501414 382454
rect 500794 382134 501414 382218
rect 500794 381898 500826 382134
rect 501062 381898 501146 382134
rect 501382 381898 501414 382134
rect 500794 342454 501414 381898
rect 500794 342218 500826 342454
rect 501062 342218 501146 342454
rect 501382 342218 501414 342454
rect 500794 342134 501414 342218
rect 500794 341898 500826 342134
rect 501062 341898 501146 342134
rect 501382 341898 501414 342134
rect 500794 302454 501414 341898
rect 500794 302218 500826 302454
rect 501062 302218 501146 302454
rect 501382 302218 501414 302454
rect 500794 302134 501414 302218
rect 500794 301898 500826 302134
rect 501062 301898 501146 302134
rect 501382 301898 501414 302134
rect 500794 262454 501414 301898
rect 500794 262218 500826 262454
rect 501062 262218 501146 262454
rect 501382 262218 501414 262454
rect 500794 262134 501414 262218
rect 500794 261898 500826 262134
rect 501062 261898 501146 262134
rect 501382 261898 501414 262134
rect 500794 222454 501414 261898
rect 500794 222218 500826 222454
rect 501062 222218 501146 222454
rect 501382 222218 501414 222454
rect 500794 222134 501414 222218
rect 500794 221898 500826 222134
rect 501062 221898 501146 222134
rect 501382 221898 501414 222134
rect 500794 182454 501414 221898
rect 500794 182218 500826 182454
rect 501062 182218 501146 182454
rect 501382 182218 501414 182454
rect 500794 182134 501414 182218
rect 500794 181898 500826 182134
rect 501062 181898 501146 182134
rect 501382 181898 501414 182134
rect 500794 142454 501414 181898
rect 500794 142218 500826 142454
rect 501062 142218 501146 142454
rect 501382 142218 501414 142454
rect 500794 142134 501414 142218
rect 500794 141898 500826 142134
rect 501062 141898 501146 142134
rect 501382 141898 501414 142134
rect 500794 102454 501414 141898
rect 500794 102218 500826 102454
rect 501062 102218 501146 102454
rect 501382 102218 501414 102454
rect 500794 102134 501414 102218
rect 500794 101898 500826 102134
rect 501062 101898 501146 102134
rect 501382 101898 501414 102134
rect 500794 62454 501414 101898
rect 500794 62218 500826 62454
rect 501062 62218 501146 62454
rect 501382 62218 501414 62454
rect 500794 62134 501414 62218
rect 500794 61898 500826 62134
rect 501062 61898 501146 62134
rect 501382 61898 501414 62134
rect 500794 22454 501414 61898
rect 500794 22218 500826 22454
rect 501062 22218 501146 22454
rect 501382 22218 501414 22454
rect 500794 22134 501414 22218
rect 500794 21898 500826 22134
rect 501062 21898 501146 22134
rect 501382 21898 501414 22134
rect 500794 -1306 501414 21898
rect 500794 -1542 500826 -1306
rect 501062 -1542 501146 -1306
rect 501382 -1542 501414 -1306
rect 500794 -1626 501414 -1542
rect 500794 -1862 500826 -1626
rect 501062 -1862 501146 -1626
rect 501382 -1862 501414 -1626
rect 500794 -1894 501414 -1862
rect 504514 666174 505134 707162
rect 504514 665938 504546 666174
rect 504782 665938 504866 666174
rect 505102 665938 505134 666174
rect 504514 665854 505134 665938
rect 504514 665618 504546 665854
rect 504782 665618 504866 665854
rect 505102 665618 505134 665854
rect 504514 626174 505134 665618
rect 504514 625938 504546 626174
rect 504782 625938 504866 626174
rect 505102 625938 505134 626174
rect 504514 625854 505134 625938
rect 504514 625618 504546 625854
rect 504782 625618 504866 625854
rect 505102 625618 505134 625854
rect 504514 586174 505134 625618
rect 504514 585938 504546 586174
rect 504782 585938 504866 586174
rect 505102 585938 505134 586174
rect 504514 585854 505134 585938
rect 504514 585618 504546 585854
rect 504782 585618 504866 585854
rect 505102 585618 505134 585854
rect 504514 546174 505134 585618
rect 504514 545938 504546 546174
rect 504782 545938 504866 546174
rect 505102 545938 505134 546174
rect 504514 545854 505134 545938
rect 504514 545618 504546 545854
rect 504782 545618 504866 545854
rect 505102 545618 505134 545854
rect 504514 506174 505134 545618
rect 504514 505938 504546 506174
rect 504782 505938 504866 506174
rect 505102 505938 505134 506174
rect 504514 505854 505134 505938
rect 504514 505618 504546 505854
rect 504782 505618 504866 505854
rect 505102 505618 505134 505854
rect 504514 466174 505134 505618
rect 504514 465938 504546 466174
rect 504782 465938 504866 466174
rect 505102 465938 505134 466174
rect 504514 465854 505134 465938
rect 504514 465618 504546 465854
rect 504782 465618 504866 465854
rect 505102 465618 505134 465854
rect 504514 426174 505134 465618
rect 504514 425938 504546 426174
rect 504782 425938 504866 426174
rect 505102 425938 505134 426174
rect 504514 425854 505134 425938
rect 504514 425618 504546 425854
rect 504782 425618 504866 425854
rect 505102 425618 505134 425854
rect 504514 386174 505134 425618
rect 504514 385938 504546 386174
rect 504782 385938 504866 386174
rect 505102 385938 505134 386174
rect 504514 385854 505134 385938
rect 504514 385618 504546 385854
rect 504782 385618 504866 385854
rect 505102 385618 505134 385854
rect 504514 346174 505134 385618
rect 504514 345938 504546 346174
rect 504782 345938 504866 346174
rect 505102 345938 505134 346174
rect 504514 345854 505134 345938
rect 504514 345618 504546 345854
rect 504782 345618 504866 345854
rect 505102 345618 505134 345854
rect 504514 306174 505134 345618
rect 504514 305938 504546 306174
rect 504782 305938 504866 306174
rect 505102 305938 505134 306174
rect 504514 305854 505134 305938
rect 504514 305618 504546 305854
rect 504782 305618 504866 305854
rect 505102 305618 505134 305854
rect 504514 266174 505134 305618
rect 504514 265938 504546 266174
rect 504782 265938 504866 266174
rect 505102 265938 505134 266174
rect 504514 265854 505134 265938
rect 504514 265618 504546 265854
rect 504782 265618 504866 265854
rect 505102 265618 505134 265854
rect 504514 226174 505134 265618
rect 504514 225938 504546 226174
rect 504782 225938 504866 226174
rect 505102 225938 505134 226174
rect 504514 225854 505134 225938
rect 504514 225618 504546 225854
rect 504782 225618 504866 225854
rect 505102 225618 505134 225854
rect 504514 186174 505134 225618
rect 504514 185938 504546 186174
rect 504782 185938 504866 186174
rect 505102 185938 505134 186174
rect 504514 185854 505134 185938
rect 504514 185618 504546 185854
rect 504782 185618 504866 185854
rect 505102 185618 505134 185854
rect 504514 146174 505134 185618
rect 504514 145938 504546 146174
rect 504782 145938 504866 146174
rect 505102 145938 505134 146174
rect 504514 145854 505134 145938
rect 504514 145618 504546 145854
rect 504782 145618 504866 145854
rect 505102 145618 505134 145854
rect 504514 106174 505134 145618
rect 504514 105938 504546 106174
rect 504782 105938 504866 106174
rect 505102 105938 505134 106174
rect 504514 105854 505134 105938
rect 504514 105618 504546 105854
rect 504782 105618 504866 105854
rect 505102 105618 505134 105854
rect 504514 66174 505134 105618
rect 504514 65938 504546 66174
rect 504782 65938 504866 66174
rect 505102 65938 505134 66174
rect 504514 65854 505134 65938
rect 504514 65618 504546 65854
rect 504782 65618 504866 65854
rect 505102 65618 505134 65854
rect 504514 26174 505134 65618
rect 504514 25938 504546 26174
rect 504782 25938 504866 26174
rect 505102 25938 505134 26174
rect 504514 25854 505134 25938
rect 504514 25618 504546 25854
rect 504782 25618 504866 25854
rect 505102 25618 505134 25854
rect 504514 -3226 505134 25618
rect 504514 -3462 504546 -3226
rect 504782 -3462 504866 -3226
rect 505102 -3462 505134 -3226
rect 504514 -3546 505134 -3462
rect 504514 -3782 504546 -3546
rect 504782 -3782 504866 -3546
rect 505102 -3782 505134 -3546
rect 504514 -3814 505134 -3782
rect 508234 669894 508854 709082
rect 508234 669658 508266 669894
rect 508502 669658 508586 669894
rect 508822 669658 508854 669894
rect 508234 669574 508854 669658
rect 508234 669338 508266 669574
rect 508502 669338 508586 669574
rect 508822 669338 508854 669574
rect 508234 629894 508854 669338
rect 508234 629658 508266 629894
rect 508502 629658 508586 629894
rect 508822 629658 508854 629894
rect 508234 629574 508854 629658
rect 508234 629338 508266 629574
rect 508502 629338 508586 629574
rect 508822 629338 508854 629574
rect 508234 589894 508854 629338
rect 508234 589658 508266 589894
rect 508502 589658 508586 589894
rect 508822 589658 508854 589894
rect 508234 589574 508854 589658
rect 508234 589338 508266 589574
rect 508502 589338 508586 589574
rect 508822 589338 508854 589574
rect 508234 549894 508854 589338
rect 508234 549658 508266 549894
rect 508502 549658 508586 549894
rect 508822 549658 508854 549894
rect 508234 549574 508854 549658
rect 508234 549338 508266 549574
rect 508502 549338 508586 549574
rect 508822 549338 508854 549574
rect 508234 509894 508854 549338
rect 508234 509658 508266 509894
rect 508502 509658 508586 509894
rect 508822 509658 508854 509894
rect 508234 509574 508854 509658
rect 508234 509338 508266 509574
rect 508502 509338 508586 509574
rect 508822 509338 508854 509574
rect 508234 469894 508854 509338
rect 508234 469658 508266 469894
rect 508502 469658 508586 469894
rect 508822 469658 508854 469894
rect 508234 469574 508854 469658
rect 508234 469338 508266 469574
rect 508502 469338 508586 469574
rect 508822 469338 508854 469574
rect 508234 429894 508854 469338
rect 508234 429658 508266 429894
rect 508502 429658 508586 429894
rect 508822 429658 508854 429894
rect 508234 429574 508854 429658
rect 508234 429338 508266 429574
rect 508502 429338 508586 429574
rect 508822 429338 508854 429574
rect 508234 389894 508854 429338
rect 508234 389658 508266 389894
rect 508502 389658 508586 389894
rect 508822 389658 508854 389894
rect 508234 389574 508854 389658
rect 508234 389338 508266 389574
rect 508502 389338 508586 389574
rect 508822 389338 508854 389574
rect 508234 349894 508854 389338
rect 508234 349658 508266 349894
rect 508502 349658 508586 349894
rect 508822 349658 508854 349894
rect 508234 349574 508854 349658
rect 508234 349338 508266 349574
rect 508502 349338 508586 349574
rect 508822 349338 508854 349574
rect 508234 309894 508854 349338
rect 508234 309658 508266 309894
rect 508502 309658 508586 309894
rect 508822 309658 508854 309894
rect 508234 309574 508854 309658
rect 508234 309338 508266 309574
rect 508502 309338 508586 309574
rect 508822 309338 508854 309574
rect 508234 269894 508854 309338
rect 508234 269658 508266 269894
rect 508502 269658 508586 269894
rect 508822 269658 508854 269894
rect 508234 269574 508854 269658
rect 508234 269338 508266 269574
rect 508502 269338 508586 269574
rect 508822 269338 508854 269574
rect 508234 229894 508854 269338
rect 508234 229658 508266 229894
rect 508502 229658 508586 229894
rect 508822 229658 508854 229894
rect 508234 229574 508854 229658
rect 508234 229338 508266 229574
rect 508502 229338 508586 229574
rect 508822 229338 508854 229574
rect 508234 189894 508854 229338
rect 508234 189658 508266 189894
rect 508502 189658 508586 189894
rect 508822 189658 508854 189894
rect 508234 189574 508854 189658
rect 508234 189338 508266 189574
rect 508502 189338 508586 189574
rect 508822 189338 508854 189574
rect 508234 149894 508854 189338
rect 508234 149658 508266 149894
rect 508502 149658 508586 149894
rect 508822 149658 508854 149894
rect 508234 149574 508854 149658
rect 508234 149338 508266 149574
rect 508502 149338 508586 149574
rect 508822 149338 508854 149574
rect 508234 109894 508854 149338
rect 508234 109658 508266 109894
rect 508502 109658 508586 109894
rect 508822 109658 508854 109894
rect 508234 109574 508854 109658
rect 508234 109338 508266 109574
rect 508502 109338 508586 109574
rect 508822 109338 508854 109574
rect 508234 69894 508854 109338
rect 508234 69658 508266 69894
rect 508502 69658 508586 69894
rect 508822 69658 508854 69894
rect 508234 69574 508854 69658
rect 508234 69338 508266 69574
rect 508502 69338 508586 69574
rect 508822 69338 508854 69574
rect 508234 29894 508854 69338
rect 508234 29658 508266 29894
rect 508502 29658 508586 29894
rect 508822 29658 508854 29894
rect 508234 29574 508854 29658
rect 508234 29338 508266 29574
rect 508502 29338 508586 29574
rect 508822 29338 508854 29574
rect 508234 -5146 508854 29338
rect 508234 -5382 508266 -5146
rect 508502 -5382 508586 -5146
rect 508822 -5382 508854 -5146
rect 508234 -5466 508854 -5382
rect 508234 -5702 508266 -5466
rect 508502 -5702 508586 -5466
rect 508822 -5702 508854 -5466
rect 508234 -5734 508854 -5702
rect 511954 673614 512574 711002
rect 531954 710598 532574 711590
rect 531954 710362 531986 710598
rect 532222 710362 532306 710598
rect 532542 710362 532574 710598
rect 531954 710278 532574 710362
rect 531954 710042 531986 710278
rect 532222 710042 532306 710278
rect 532542 710042 532574 710278
rect 528234 708678 528854 709670
rect 528234 708442 528266 708678
rect 528502 708442 528586 708678
rect 528822 708442 528854 708678
rect 528234 708358 528854 708442
rect 528234 708122 528266 708358
rect 528502 708122 528586 708358
rect 528822 708122 528854 708358
rect 524514 706758 525134 707750
rect 524514 706522 524546 706758
rect 524782 706522 524866 706758
rect 525102 706522 525134 706758
rect 524514 706438 525134 706522
rect 524514 706202 524546 706438
rect 524782 706202 524866 706438
rect 525102 706202 525134 706438
rect 511954 673378 511986 673614
rect 512222 673378 512306 673614
rect 512542 673378 512574 673614
rect 511954 673294 512574 673378
rect 511954 673058 511986 673294
rect 512222 673058 512306 673294
rect 512542 673058 512574 673294
rect 511954 633614 512574 673058
rect 511954 633378 511986 633614
rect 512222 633378 512306 633614
rect 512542 633378 512574 633614
rect 511954 633294 512574 633378
rect 511954 633058 511986 633294
rect 512222 633058 512306 633294
rect 512542 633058 512574 633294
rect 511954 593614 512574 633058
rect 511954 593378 511986 593614
rect 512222 593378 512306 593614
rect 512542 593378 512574 593614
rect 511954 593294 512574 593378
rect 511954 593058 511986 593294
rect 512222 593058 512306 593294
rect 512542 593058 512574 593294
rect 511954 553614 512574 593058
rect 511954 553378 511986 553614
rect 512222 553378 512306 553614
rect 512542 553378 512574 553614
rect 511954 553294 512574 553378
rect 511954 553058 511986 553294
rect 512222 553058 512306 553294
rect 512542 553058 512574 553294
rect 511954 513614 512574 553058
rect 511954 513378 511986 513614
rect 512222 513378 512306 513614
rect 512542 513378 512574 513614
rect 511954 513294 512574 513378
rect 511954 513058 511986 513294
rect 512222 513058 512306 513294
rect 512542 513058 512574 513294
rect 511954 473614 512574 513058
rect 511954 473378 511986 473614
rect 512222 473378 512306 473614
rect 512542 473378 512574 473614
rect 511954 473294 512574 473378
rect 511954 473058 511986 473294
rect 512222 473058 512306 473294
rect 512542 473058 512574 473294
rect 511954 433614 512574 473058
rect 511954 433378 511986 433614
rect 512222 433378 512306 433614
rect 512542 433378 512574 433614
rect 511954 433294 512574 433378
rect 511954 433058 511986 433294
rect 512222 433058 512306 433294
rect 512542 433058 512574 433294
rect 511954 393614 512574 433058
rect 511954 393378 511986 393614
rect 512222 393378 512306 393614
rect 512542 393378 512574 393614
rect 511954 393294 512574 393378
rect 511954 393058 511986 393294
rect 512222 393058 512306 393294
rect 512542 393058 512574 393294
rect 511954 353614 512574 393058
rect 511954 353378 511986 353614
rect 512222 353378 512306 353614
rect 512542 353378 512574 353614
rect 511954 353294 512574 353378
rect 511954 353058 511986 353294
rect 512222 353058 512306 353294
rect 512542 353058 512574 353294
rect 511954 313614 512574 353058
rect 511954 313378 511986 313614
rect 512222 313378 512306 313614
rect 512542 313378 512574 313614
rect 511954 313294 512574 313378
rect 511954 313058 511986 313294
rect 512222 313058 512306 313294
rect 512542 313058 512574 313294
rect 511954 273614 512574 313058
rect 511954 273378 511986 273614
rect 512222 273378 512306 273614
rect 512542 273378 512574 273614
rect 511954 273294 512574 273378
rect 511954 273058 511986 273294
rect 512222 273058 512306 273294
rect 512542 273058 512574 273294
rect 511954 233614 512574 273058
rect 511954 233378 511986 233614
rect 512222 233378 512306 233614
rect 512542 233378 512574 233614
rect 511954 233294 512574 233378
rect 511954 233058 511986 233294
rect 512222 233058 512306 233294
rect 512542 233058 512574 233294
rect 511954 193614 512574 233058
rect 511954 193378 511986 193614
rect 512222 193378 512306 193614
rect 512542 193378 512574 193614
rect 511954 193294 512574 193378
rect 511954 193058 511986 193294
rect 512222 193058 512306 193294
rect 512542 193058 512574 193294
rect 511954 153614 512574 193058
rect 511954 153378 511986 153614
rect 512222 153378 512306 153614
rect 512542 153378 512574 153614
rect 511954 153294 512574 153378
rect 511954 153058 511986 153294
rect 512222 153058 512306 153294
rect 512542 153058 512574 153294
rect 511954 113614 512574 153058
rect 511954 113378 511986 113614
rect 512222 113378 512306 113614
rect 512542 113378 512574 113614
rect 511954 113294 512574 113378
rect 511954 113058 511986 113294
rect 512222 113058 512306 113294
rect 512542 113058 512574 113294
rect 511954 73614 512574 113058
rect 511954 73378 511986 73614
rect 512222 73378 512306 73614
rect 512542 73378 512574 73614
rect 511954 73294 512574 73378
rect 511954 73058 511986 73294
rect 512222 73058 512306 73294
rect 512542 73058 512574 73294
rect 511954 33614 512574 73058
rect 511954 33378 511986 33614
rect 512222 33378 512306 33614
rect 512542 33378 512574 33614
rect 511954 33294 512574 33378
rect 511954 33058 511986 33294
rect 512222 33058 512306 33294
rect 512542 33058 512574 33294
rect 491954 -6342 491986 -6106
rect 492222 -6342 492306 -6106
rect 492542 -6342 492574 -6106
rect 491954 -6426 492574 -6342
rect 491954 -6662 491986 -6426
rect 492222 -6662 492306 -6426
rect 492542 -6662 492574 -6426
rect 491954 -7654 492574 -6662
rect 511954 -7066 512574 33058
rect 520794 704838 521414 705830
rect 520794 704602 520826 704838
rect 521062 704602 521146 704838
rect 521382 704602 521414 704838
rect 520794 704518 521414 704602
rect 520794 704282 520826 704518
rect 521062 704282 521146 704518
rect 521382 704282 521414 704518
rect 520794 682454 521414 704282
rect 520794 682218 520826 682454
rect 521062 682218 521146 682454
rect 521382 682218 521414 682454
rect 520794 682134 521414 682218
rect 520794 681898 520826 682134
rect 521062 681898 521146 682134
rect 521382 681898 521414 682134
rect 520794 642454 521414 681898
rect 520794 642218 520826 642454
rect 521062 642218 521146 642454
rect 521382 642218 521414 642454
rect 520794 642134 521414 642218
rect 520794 641898 520826 642134
rect 521062 641898 521146 642134
rect 521382 641898 521414 642134
rect 520794 602454 521414 641898
rect 520794 602218 520826 602454
rect 521062 602218 521146 602454
rect 521382 602218 521414 602454
rect 520794 602134 521414 602218
rect 520794 601898 520826 602134
rect 521062 601898 521146 602134
rect 521382 601898 521414 602134
rect 520794 562454 521414 601898
rect 520794 562218 520826 562454
rect 521062 562218 521146 562454
rect 521382 562218 521414 562454
rect 520794 562134 521414 562218
rect 520794 561898 520826 562134
rect 521062 561898 521146 562134
rect 521382 561898 521414 562134
rect 520794 522454 521414 561898
rect 520794 522218 520826 522454
rect 521062 522218 521146 522454
rect 521382 522218 521414 522454
rect 520794 522134 521414 522218
rect 520794 521898 520826 522134
rect 521062 521898 521146 522134
rect 521382 521898 521414 522134
rect 520794 482454 521414 521898
rect 520794 482218 520826 482454
rect 521062 482218 521146 482454
rect 521382 482218 521414 482454
rect 520794 482134 521414 482218
rect 520794 481898 520826 482134
rect 521062 481898 521146 482134
rect 521382 481898 521414 482134
rect 520794 442454 521414 481898
rect 520794 442218 520826 442454
rect 521062 442218 521146 442454
rect 521382 442218 521414 442454
rect 520794 442134 521414 442218
rect 520794 441898 520826 442134
rect 521062 441898 521146 442134
rect 521382 441898 521414 442134
rect 520794 402454 521414 441898
rect 520794 402218 520826 402454
rect 521062 402218 521146 402454
rect 521382 402218 521414 402454
rect 520794 402134 521414 402218
rect 520794 401898 520826 402134
rect 521062 401898 521146 402134
rect 521382 401898 521414 402134
rect 520794 362454 521414 401898
rect 520794 362218 520826 362454
rect 521062 362218 521146 362454
rect 521382 362218 521414 362454
rect 520794 362134 521414 362218
rect 520794 361898 520826 362134
rect 521062 361898 521146 362134
rect 521382 361898 521414 362134
rect 520794 322454 521414 361898
rect 520794 322218 520826 322454
rect 521062 322218 521146 322454
rect 521382 322218 521414 322454
rect 520794 322134 521414 322218
rect 520794 321898 520826 322134
rect 521062 321898 521146 322134
rect 521382 321898 521414 322134
rect 520794 282454 521414 321898
rect 520794 282218 520826 282454
rect 521062 282218 521146 282454
rect 521382 282218 521414 282454
rect 520794 282134 521414 282218
rect 520794 281898 520826 282134
rect 521062 281898 521146 282134
rect 521382 281898 521414 282134
rect 520794 242454 521414 281898
rect 520794 242218 520826 242454
rect 521062 242218 521146 242454
rect 521382 242218 521414 242454
rect 520794 242134 521414 242218
rect 520794 241898 520826 242134
rect 521062 241898 521146 242134
rect 521382 241898 521414 242134
rect 520794 202454 521414 241898
rect 520794 202218 520826 202454
rect 521062 202218 521146 202454
rect 521382 202218 521414 202454
rect 520794 202134 521414 202218
rect 520794 201898 520826 202134
rect 521062 201898 521146 202134
rect 521382 201898 521414 202134
rect 520794 162454 521414 201898
rect 520794 162218 520826 162454
rect 521062 162218 521146 162454
rect 521382 162218 521414 162454
rect 520794 162134 521414 162218
rect 520794 161898 520826 162134
rect 521062 161898 521146 162134
rect 521382 161898 521414 162134
rect 520794 122454 521414 161898
rect 520794 122218 520826 122454
rect 521062 122218 521146 122454
rect 521382 122218 521414 122454
rect 520794 122134 521414 122218
rect 520794 121898 520826 122134
rect 521062 121898 521146 122134
rect 521382 121898 521414 122134
rect 520794 82454 521414 121898
rect 520794 82218 520826 82454
rect 521062 82218 521146 82454
rect 521382 82218 521414 82454
rect 520794 82134 521414 82218
rect 520794 81898 520826 82134
rect 521062 81898 521146 82134
rect 521382 81898 521414 82134
rect 520794 42454 521414 81898
rect 520794 42218 520826 42454
rect 521062 42218 521146 42454
rect 521382 42218 521414 42454
rect 520794 42134 521414 42218
rect 520794 41898 520826 42134
rect 521062 41898 521146 42134
rect 521382 41898 521414 42134
rect 520794 2454 521414 41898
rect 520794 2218 520826 2454
rect 521062 2218 521146 2454
rect 521382 2218 521414 2454
rect 520794 2134 521414 2218
rect 520794 1898 520826 2134
rect 521062 1898 521146 2134
rect 521382 1898 521414 2134
rect 520794 -346 521414 1898
rect 520794 -582 520826 -346
rect 521062 -582 521146 -346
rect 521382 -582 521414 -346
rect 520794 -666 521414 -582
rect 520794 -902 520826 -666
rect 521062 -902 521146 -666
rect 521382 -902 521414 -666
rect 520794 -1894 521414 -902
rect 524514 686174 525134 706202
rect 524514 685938 524546 686174
rect 524782 685938 524866 686174
rect 525102 685938 525134 686174
rect 524514 685854 525134 685938
rect 524514 685618 524546 685854
rect 524782 685618 524866 685854
rect 525102 685618 525134 685854
rect 524514 646174 525134 685618
rect 524514 645938 524546 646174
rect 524782 645938 524866 646174
rect 525102 645938 525134 646174
rect 524514 645854 525134 645938
rect 524514 645618 524546 645854
rect 524782 645618 524866 645854
rect 525102 645618 525134 645854
rect 524514 606174 525134 645618
rect 524514 605938 524546 606174
rect 524782 605938 524866 606174
rect 525102 605938 525134 606174
rect 524514 605854 525134 605938
rect 524514 605618 524546 605854
rect 524782 605618 524866 605854
rect 525102 605618 525134 605854
rect 524514 566174 525134 605618
rect 524514 565938 524546 566174
rect 524782 565938 524866 566174
rect 525102 565938 525134 566174
rect 524514 565854 525134 565938
rect 524514 565618 524546 565854
rect 524782 565618 524866 565854
rect 525102 565618 525134 565854
rect 524514 526174 525134 565618
rect 524514 525938 524546 526174
rect 524782 525938 524866 526174
rect 525102 525938 525134 526174
rect 524514 525854 525134 525938
rect 524514 525618 524546 525854
rect 524782 525618 524866 525854
rect 525102 525618 525134 525854
rect 524514 486174 525134 525618
rect 524514 485938 524546 486174
rect 524782 485938 524866 486174
rect 525102 485938 525134 486174
rect 524514 485854 525134 485938
rect 524514 485618 524546 485854
rect 524782 485618 524866 485854
rect 525102 485618 525134 485854
rect 524514 446174 525134 485618
rect 524514 445938 524546 446174
rect 524782 445938 524866 446174
rect 525102 445938 525134 446174
rect 524514 445854 525134 445938
rect 524514 445618 524546 445854
rect 524782 445618 524866 445854
rect 525102 445618 525134 445854
rect 524514 406174 525134 445618
rect 524514 405938 524546 406174
rect 524782 405938 524866 406174
rect 525102 405938 525134 406174
rect 524514 405854 525134 405938
rect 524514 405618 524546 405854
rect 524782 405618 524866 405854
rect 525102 405618 525134 405854
rect 524514 366174 525134 405618
rect 524514 365938 524546 366174
rect 524782 365938 524866 366174
rect 525102 365938 525134 366174
rect 524514 365854 525134 365938
rect 524514 365618 524546 365854
rect 524782 365618 524866 365854
rect 525102 365618 525134 365854
rect 524514 326174 525134 365618
rect 524514 325938 524546 326174
rect 524782 325938 524866 326174
rect 525102 325938 525134 326174
rect 524514 325854 525134 325938
rect 524514 325618 524546 325854
rect 524782 325618 524866 325854
rect 525102 325618 525134 325854
rect 524514 286174 525134 325618
rect 524514 285938 524546 286174
rect 524782 285938 524866 286174
rect 525102 285938 525134 286174
rect 524514 285854 525134 285938
rect 524514 285618 524546 285854
rect 524782 285618 524866 285854
rect 525102 285618 525134 285854
rect 524514 246174 525134 285618
rect 524514 245938 524546 246174
rect 524782 245938 524866 246174
rect 525102 245938 525134 246174
rect 524514 245854 525134 245938
rect 524514 245618 524546 245854
rect 524782 245618 524866 245854
rect 525102 245618 525134 245854
rect 524514 206174 525134 245618
rect 524514 205938 524546 206174
rect 524782 205938 524866 206174
rect 525102 205938 525134 206174
rect 524514 205854 525134 205938
rect 524514 205618 524546 205854
rect 524782 205618 524866 205854
rect 525102 205618 525134 205854
rect 524514 166174 525134 205618
rect 524514 165938 524546 166174
rect 524782 165938 524866 166174
rect 525102 165938 525134 166174
rect 524514 165854 525134 165938
rect 524514 165618 524546 165854
rect 524782 165618 524866 165854
rect 525102 165618 525134 165854
rect 524514 126174 525134 165618
rect 524514 125938 524546 126174
rect 524782 125938 524866 126174
rect 525102 125938 525134 126174
rect 524514 125854 525134 125938
rect 524514 125618 524546 125854
rect 524782 125618 524866 125854
rect 525102 125618 525134 125854
rect 524514 86174 525134 125618
rect 524514 85938 524546 86174
rect 524782 85938 524866 86174
rect 525102 85938 525134 86174
rect 524514 85854 525134 85938
rect 524514 85618 524546 85854
rect 524782 85618 524866 85854
rect 525102 85618 525134 85854
rect 524514 46174 525134 85618
rect 524514 45938 524546 46174
rect 524782 45938 524866 46174
rect 525102 45938 525134 46174
rect 524514 45854 525134 45938
rect 524514 45618 524546 45854
rect 524782 45618 524866 45854
rect 525102 45618 525134 45854
rect 524514 6174 525134 45618
rect 524514 5938 524546 6174
rect 524782 5938 524866 6174
rect 525102 5938 525134 6174
rect 524514 5854 525134 5938
rect 524514 5618 524546 5854
rect 524782 5618 524866 5854
rect 525102 5618 525134 5854
rect 524514 -2266 525134 5618
rect 524514 -2502 524546 -2266
rect 524782 -2502 524866 -2266
rect 525102 -2502 525134 -2266
rect 524514 -2586 525134 -2502
rect 524514 -2822 524546 -2586
rect 524782 -2822 524866 -2586
rect 525102 -2822 525134 -2586
rect 524514 -3814 525134 -2822
rect 528234 689894 528854 708122
rect 528234 689658 528266 689894
rect 528502 689658 528586 689894
rect 528822 689658 528854 689894
rect 528234 689574 528854 689658
rect 528234 689338 528266 689574
rect 528502 689338 528586 689574
rect 528822 689338 528854 689574
rect 528234 649894 528854 689338
rect 528234 649658 528266 649894
rect 528502 649658 528586 649894
rect 528822 649658 528854 649894
rect 528234 649574 528854 649658
rect 528234 649338 528266 649574
rect 528502 649338 528586 649574
rect 528822 649338 528854 649574
rect 528234 609894 528854 649338
rect 528234 609658 528266 609894
rect 528502 609658 528586 609894
rect 528822 609658 528854 609894
rect 528234 609574 528854 609658
rect 528234 609338 528266 609574
rect 528502 609338 528586 609574
rect 528822 609338 528854 609574
rect 528234 569894 528854 609338
rect 528234 569658 528266 569894
rect 528502 569658 528586 569894
rect 528822 569658 528854 569894
rect 528234 569574 528854 569658
rect 528234 569338 528266 569574
rect 528502 569338 528586 569574
rect 528822 569338 528854 569574
rect 528234 529894 528854 569338
rect 528234 529658 528266 529894
rect 528502 529658 528586 529894
rect 528822 529658 528854 529894
rect 528234 529574 528854 529658
rect 528234 529338 528266 529574
rect 528502 529338 528586 529574
rect 528822 529338 528854 529574
rect 528234 489894 528854 529338
rect 528234 489658 528266 489894
rect 528502 489658 528586 489894
rect 528822 489658 528854 489894
rect 528234 489574 528854 489658
rect 528234 489338 528266 489574
rect 528502 489338 528586 489574
rect 528822 489338 528854 489574
rect 528234 449894 528854 489338
rect 528234 449658 528266 449894
rect 528502 449658 528586 449894
rect 528822 449658 528854 449894
rect 528234 449574 528854 449658
rect 528234 449338 528266 449574
rect 528502 449338 528586 449574
rect 528822 449338 528854 449574
rect 528234 409894 528854 449338
rect 528234 409658 528266 409894
rect 528502 409658 528586 409894
rect 528822 409658 528854 409894
rect 528234 409574 528854 409658
rect 528234 409338 528266 409574
rect 528502 409338 528586 409574
rect 528822 409338 528854 409574
rect 528234 369894 528854 409338
rect 528234 369658 528266 369894
rect 528502 369658 528586 369894
rect 528822 369658 528854 369894
rect 528234 369574 528854 369658
rect 528234 369338 528266 369574
rect 528502 369338 528586 369574
rect 528822 369338 528854 369574
rect 528234 329894 528854 369338
rect 528234 329658 528266 329894
rect 528502 329658 528586 329894
rect 528822 329658 528854 329894
rect 528234 329574 528854 329658
rect 528234 329338 528266 329574
rect 528502 329338 528586 329574
rect 528822 329338 528854 329574
rect 528234 289894 528854 329338
rect 528234 289658 528266 289894
rect 528502 289658 528586 289894
rect 528822 289658 528854 289894
rect 528234 289574 528854 289658
rect 528234 289338 528266 289574
rect 528502 289338 528586 289574
rect 528822 289338 528854 289574
rect 528234 249894 528854 289338
rect 528234 249658 528266 249894
rect 528502 249658 528586 249894
rect 528822 249658 528854 249894
rect 528234 249574 528854 249658
rect 528234 249338 528266 249574
rect 528502 249338 528586 249574
rect 528822 249338 528854 249574
rect 528234 209894 528854 249338
rect 528234 209658 528266 209894
rect 528502 209658 528586 209894
rect 528822 209658 528854 209894
rect 528234 209574 528854 209658
rect 528234 209338 528266 209574
rect 528502 209338 528586 209574
rect 528822 209338 528854 209574
rect 528234 169894 528854 209338
rect 528234 169658 528266 169894
rect 528502 169658 528586 169894
rect 528822 169658 528854 169894
rect 528234 169574 528854 169658
rect 528234 169338 528266 169574
rect 528502 169338 528586 169574
rect 528822 169338 528854 169574
rect 528234 129894 528854 169338
rect 528234 129658 528266 129894
rect 528502 129658 528586 129894
rect 528822 129658 528854 129894
rect 528234 129574 528854 129658
rect 528234 129338 528266 129574
rect 528502 129338 528586 129574
rect 528822 129338 528854 129574
rect 528234 89894 528854 129338
rect 528234 89658 528266 89894
rect 528502 89658 528586 89894
rect 528822 89658 528854 89894
rect 528234 89574 528854 89658
rect 528234 89338 528266 89574
rect 528502 89338 528586 89574
rect 528822 89338 528854 89574
rect 528234 49894 528854 89338
rect 528234 49658 528266 49894
rect 528502 49658 528586 49894
rect 528822 49658 528854 49894
rect 528234 49574 528854 49658
rect 528234 49338 528266 49574
rect 528502 49338 528586 49574
rect 528822 49338 528854 49574
rect 528234 9894 528854 49338
rect 528234 9658 528266 9894
rect 528502 9658 528586 9894
rect 528822 9658 528854 9894
rect 528234 9574 528854 9658
rect 528234 9338 528266 9574
rect 528502 9338 528586 9574
rect 528822 9338 528854 9574
rect 528234 -4186 528854 9338
rect 528234 -4422 528266 -4186
rect 528502 -4422 528586 -4186
rect 528822 -4422 528854 -4186
rect 528234 -4506 528854 -4422
rect 528234 -4742 528266 -4506
rect 528502 -4742 528586 -4506
rect 528822 -4742 528854 -4506
rect 528234 -5734 528854 -4742
rect 531954 693614 532574 710042
rect 551954 711558 552574 711590
rect 551954 711322 551986 711558
rect 552222 711322 552306 711558
rect 552542 711322 552574 711558
rect 551954 711238 552574 711322
rect 551954 711002 551986 711238
rect 552222 711002 552306 711238
rect 552542 711002 552574 711238
rect 548234 709638 548854 709670
rect 548234 709402 548266 709638
rect 548502 709402 548586 709638
rect 548822 709402 548854 709638
rect 548234 709318 548854 709402
rect 548234 709082 548266 709318
rect 548502 709082 548586 709318
rect 548822 709082 548854 709318
rect 544514 707718 545134 707750
rect 544514 707482 544546 707718
rect 544782 707482 544866 707718
rect 545102 707482 545134 707718
rect 544514 707398 545134 707482
rect 544514 707162 544546 707398
rect 544782 707162 544866 707398
rect 545102 707162 545134 707398
rect 531954 693378 531986 693614
rect 532222 693378 532306 693614
rect 532542 693378 532574 693614
rect 531954 693294 532574 693378
rect 531954 693058 531986 693294
rect 532222 693058 532306 693294
rect 532542 693058 532574 693294
rect 531954 653614 532574 693058
rect 531954 653378 531986 653614
rect 532222 653378 532306 653614
rect 532542 653378 532574 653614
rect 531954 653294 532574 653378
rect 531954 653058 531986 653294
rect 532222 653058 532306 653294
rect 532542 653058 532574 653294
rect 531954 613614 532574 653058
rect 531954 613378 531986 613614
rect 532222 613378 532306 613614
rect 532542 613378 532574 613614
rect 531954 613294 532574 613378
rect 531954 613058 531986 613294
rect 532222 613058 532306 613294
rect 532542 613058 532574 613294
rect 531954 573614 532574 613058
rect 531954 573378 531986 573614
rect 532222 573378 532306 573614
rect 532542 573378 532574 573614
rect 531954 573294 532574 573378
rect 531954 573058 531986 573294
rect 532222 573058 532306 573294
rect 532542 573058 532574 573294
rect 531954 533614 532574 573058
rect 531954 533378 531986 533614
rect 532222 533378 532306 533614
rect 532542 533378 532574 533614
rect 531954 533294 532574 533378
rect 531954 533058 531986 533294
rect 532222 533058 532306 533294
rect 532542 533058 532574 533294
rect 531954 493614 532574 533058
rect 531954 493378 531986 493614
rect 532222 493378 532306 493614
rect 532542 493378 532574 493614
rect 531954 493294 532574 493378
rect 531954 493058 531986 493294
rect 532222 493058 532306 493294
rect 532542 493058 532574 493294
rect 531954 453614 532574 493058
rect 531954 453378 531986 453614
rect 532222 453378 532306 453614
rect 532542 453378 532574 453614
rect 531954 453294 532574 453378
rect 531954 453058 531986 453294
rect 532222 453058 532306 453294
rect 532542 453058 532574 453294
rect 531954 413614 532574 453058
rect 531954 413378 531986 413614
rect 532222 413378 532306 413614
rect 532542 413378 532574 413614
rect 531954 413294 532574 413378
rect 531954 413058 531986 413294
rect 532222 413058 532306 413294
rect 532542 413058 532574 413294
rect 531954 373614 532574 413058
rect 531954 373378 531986 373614
rect 532222 373378 532306 373614
rect 532542 373378 532574 373614
rect 531954 373294 532574 373378
rect 531954 373058 531986 373294
rect 532222 373058 532306 373294
rect 532542 373058 532574 373294
rect 531954 333614 532574 373058
rect 531954 333378 531986 333614
rect 532222 333378 532306 333614
rect 532542 333378 532574 333614
rect 531954 333294 532574 333378
rect 531954 333058 531986 333294
rect 532222 333058 532306 333294
rect 532542 333058 532574 333294
rect 531954 293614 532574 333058
rect 531954 293378 531986 293614
rect 532222 293378 532306 293614
rect 532542 293378 532574 293614
rect 531954 293294 532574 293378
rect 531954 293058 531986 293294
rect 532222 293058 532306 293294
rect 532542 293058 532574 293294
rect 531954 253614 532574 293058
rect 531954 253378 531986 253614
rect 532222 253378 532306 253614
rect 532542 253378 532574 253614
rect 531954 253294 532574 253378
rect 531954 253058 531986 253294
rect 532222 253058 532306 253294
rect 532542 253058 532574 253294
rect 531954 213614 532574 253058
rect 531954 213378 531986 213614
rect 532222 213378 532306 213614
rect 532542 213378 532574 213614
rect 531954 213294 532574 213378
rect 531954 213058 531986 213294
rect 532222 213058 532306 213294
rect 532542 213058 532574 213294
rect 531954 173614 532574 213058
rect 531954 173378 531986 173614
rect 532222 173378 532306 173614
rect 532542 173378 532574 173614
rect 531954 173294 532574 173378
rect 531954 173058 531986 173294
rect 532222 173058 532306 173294
rect 532542 173058 532574 173294
rect 531954 133614 532574 173058
rect 531954 133378 531986 133614
rect 532222 133378 532306 133614
rect 532542 133378 532574 133614
rect 531954 133294 532574 133378
rect 531954 133058 531986 133294
rect 532222 133058 532306 133294
rect 532542 133058 532574 133294
rect 531954 93614 532574 133058
rect 531954 93378 531986 93614
rect 532222 93378 532306 93614
rect 532542 93378 532574 93614
rect 531954 93294 532574 93378
rect 531954 93058 531986 93294
rect 532222 93058 532306 93294
rect 532542 93058 532574 93294
rect 531954 53614 532574 93058
rect 531954 53378 531986 53614
rect 532222 53378 532306 53614
rect 532542 53378 532574 53614
rect 531954 53294 532574 53378
rect 531954 53058 531986 53294
rect 532222 53058 532306 53294
rect 532542 53058 532574 53294
rect 531954 13614 532574 53058
rect 531954 13378 531986 13614
rect 532222 13378 532306 13614
rect 532542 13378 532574 13614
rect 531954 13294 532574 13378
rect 531954 13058 531986 13294
rect 532222 13058 532306 13294
rect 532542 13058 532574 13294
rect 511954 -7302 511986 -7066
rect 512222 -7302 512306 -7066
rect 512542 -7302 512574 -7066
rect 511954 -7386 512574 -7302
rect 511954 -7622 511986 -7386
rect 512222 -7622 512306 -7386
rect 512542 -7622 512574 -7386
rect 511954 -7654 512574 -7622
rect 531954 -6106 532574 13058
rect 540794 705798 541414 705830
rect 540794 705562 540826 705798
rect 541062 705562 541146 705798
rect 541382 705562 541414 705798
rect 540794 705478 541414 705562
rect 540794 705242 540826 705478
rect 541062 705242 541146 705478
rect 541382 705242 541414 705478
rect 540794 662454 541414 705242
rect 540794 662218 540826 662454
rect 541062 662218 541146 662454
rect 541382 662218 541414 662454
rect 540794 662134 541414 662218
rect 540794 661898 540826 662134
rect 541062 661898 541146 662134
rect 541382 661898 541414 662134
rect 540794 622454 541414 661898
rect 540794 622218 540826 622454
rect 541062 622218 541146 622454
rect 541382 622218 541414 622454
rect 540794 622134 541414 622218
rect 540794 621898 540826 622134
rect 541062 621898 541146 622134
rect 541382 621898 541414 622134
rect 540794 582454 541414 621898
rect 540794 582218 540826 582454
rect 541062 582218 541146 582454
rect 541382 582218 541414 582454
rect 540794 582134 541414 582218
rect 540794 581898 540826 582134
rect 541062 581898 541146 582134
rect 541382 581898 541414 582134
rect 540794 542454 541414 581898
rect 540794 542218 540826 542454
rect 541062 542218 541146 542454
rect 541382 542218 541414 542454
rect 540794 542134 541414 542218
rect 540794 541898 540826 542134
rect 541062 541898 541146 542134
rect 541382 541898 541414 542134
rect 540794 502454 541414 541898
rect 540794 502218 540826 502454
rect 541062 502218 541146 502454
rect 541382 502218 541414 502454
rect 540794 502134 541414 502218
rect 540794 501898 540826 502134
rect 541062 501898 541146 502134
rect 541382 501898 541414 502134
rect 540794 462454 541414 501898
rect 540794 462218 540826 462454
rect 541062 462218 541146 462454
rect 541382 462218 541414 462454
rect 540794 462134 541414 462218
rect 540794 461898 540826 462134
rect 541062 461898 541146 462134
rect 541382 461898 541414 462134
rect 540794 422454 541414 461898
rect 540794 422218 540826 422454
rect 541062 422218 541146 422454
rect 541382 422218 541414 422454
rect 540794 422134 541414 422218
rect 540794 421898 540826 422134
rect 541062 421898 541146 422134
rect 541382 421898 541414 422134
rect 540794 382454 541414 421898
rect 540794 382218 540826 382454
rect 541062 382218 541146 382454
rect 541382 382218 541414 382454
rect 540794 382134 541414 382218
rect 540794 381898 540826 382134
rect 541062 381898 541146 382134
rect 541382 381898 541414 382134
rect 540794 342454 541414 381898
rect 540794 342218 540826 342454
rect 541062 342218 541146 342454
rect 541382 342218 541414 342454
rect 540794 342134 541414 342218
rect 540794 341898 540826 342134
rect 541062 341898 541146 342134
rect 541382 341898 541414 342134
rect 540794 302454 541414 341898
rect 540794 302218 540826 302454
rect 541062 302218 541146 302454
rect 541382 302218 541414 302454
rect 540794 302134 541414 302218
rect 540794 301898 540826 302134
rect 541062 301898 541146 302134
rect 541382 301898 541414 302134
rect 540794 262454 541414 301898
rect 540794 262218 540826 262454
rect 541062 262218 541146 262454
rect 541382 262218 541414 262454
rect 540794 262134 541414 262218
rect 540794 261898 540826 262134
rect 541062 261898 541146 262134
rect 541382 261898 541414 262134
rect 540794 222454 541414 261898
rect 540794 222218 540826 222454
rect 541062 222218 541146 222454
rect 541382 222218 541414 222454
rect 540794 222134 541414 222218
rect 540794 221898 540826 222134
rect 541062 221898 541146 222134
rect 541382 221898 541414 222134
rect 540794 182454 541414 221898
rect 540794 182218 540826 182454
rect 541062 182218 541146 182454
rect 541382 182218 541414 182454
rect 540794 182134 541414 182218
rect 540794 181898 540826 182134
rect 541062 181898 541146 182134
rect 541382 181898 541414 182134
rect 540794 142454 541414 181898
rect 540794 142218 540826 142454
rect 541062 142218 541146 142454
rect 541382 142218 541414 142454
rect 540794 142134 541414 142218
rect 540794 141898 540826 142134
rect 541062 141898 541146 142134
rect 541382 141898 541414 142134
rect 540794 102454 541414 141898
rect 540794 102218 540826 102454
rect 541062 102218 541146 102454
rect 541382 102218 541414 102454
rect 540794 102134 541414 102218
rect 540794 101898 540826 102134
rect 541062 101898 541146 102134
rect 541382 101898 541414 102134
rect 540794 62454 541414 101898
rect 540794 62218 540826 62454
rect 541062 62218 541146 62454
rect 541382 62218 541414 62454
rect 540794 62134 541414 62218
rect 540794 61898 540826 62134
rect 541062 61898 541146 62134
rect 541382 61898 541414 62134
rect 540794 22454 541414 61898
rect 540794 22218 540826 22454
rect 541062 22218 541146 22454
rect 541382 22218 541414 22454
rect 540794 22134 541414 22218
rect 540794 21898 540826 22134
rect 541062 21898 541146 22134
rect 541382 21898 541414 22134
rect 540794 -1306 541414 21898
rect 540794 -1542 540826 -1306
rect 541062 -1542 541146 -1306
rect 541382 -1542 541414 -1306
rect 540794 -1626 541414 -1542
rect 540794 -1862 540826 -1626
rect 541062 -1862 541146 -1626
rect 541382 -1862 541414 -1626
rect 540794 -1894 541414 -1862
rect 544514 666174 545134 707162
rect 544514 665938 544546 666174
rect 544782 665938 544866 666174
rect 545102 665938 545134 666174
rect 544514 665854 545134 665938
rect 544514 665618 544546 665854
rect 544782 665618 544866 665854
rect 545102 665618 545134 665854
rect 544514 626174 545134 665618
rect 544514 625938 544546 626174
rect 544782 625938 544866 626174
rect 545102 625938 545134 626174
rect 544514 625854 545134 625938
rect 544514 625618 544546 625854
rect 544782 625618 544866 625854
rect 545102 625618 545134 625854
rect 544514 586174 545134 625618
rect 544514 585938 544546 586174
rect 544782 585938 544866 586174
rect 545102 585938 545134 586174
rect 544514 585854 545134 585938
rect 544514 585618 544546 585854
rect 544782 585618 544866 585854
rect 545102 585618 545134 585854
rect 544514 546174 545134 585618
rect 544514 545938 544546 546174
rect 544782 545938 544866 546174
rect 545102 545938 545134 546174
rect 544514 545854 545134 545938
rect 544514 545618 544546 545854
rect 544782 545618 544866 545854
rect 545102 545618 545134 545854
rect 544514 506174 545134 545618
rect 544514 505938 544546 506174
rect 544782 505938 544866 506174
rect 545102 505938 545134 506174
rect 544514 505854 545134 505938
rect 544514 505618 544546 505854
rect 544782 505618 544866 505854
rect 545102 505618 545134 505854
rect 544514 466174 545134 505618
rect 544514 465938 544546 466174
rect 544782 465938 544866 466174
rect 545102 465938 545134 466174
rect 544514 465854 545134 465938
rect 544514 465618 544546 465854
rect 544782 465618 544866 465854
rect 545102 465618 545134 465854
rect 544514 426174 545134 465618
rect 544514 425938 544546 426174
rect 544782 425938 544866 426174
rect 545102 425938 545134 426174
rect 544514 425854 545134 425938
rect 544514 425618 544546 425854
rect 544782 425618 544866 425854
rect 545102 425618 545134 425854
rect 544514 386174 545134 425618
rect 544514 385938 544546 386174
rect 544782 385938 544866 386174
rect 545102 385938 545134 386174
rect 544514 385854 545134 385938
rect 544514 385618 544546 385854
rect 544782 385618 544866 385854
rect 545102 385618 545134 385854
rect 544514 346174 545134 385618
rect 544514 345938 544546 346174
rect 544782 345938 544866 346174
rect 545102 345938 545134 346174
rect 544514 345854 545134 345938
rect 544514 345618 544546 345854
rect 544782 345618 544866 345854
rect 545102 345618 545134 345854
rect 544514 306174 545134 345618
rect 544514 305938 544546 306174
rect 544782 305938 544866 306174
rect 545102 305938 545134 306174
rect 544514 305854 545134 305938
rect 544514 305618 544546 305854
rect 544782 305618 544866 305854
rect 545102 305618 545134 305854
rect 544514 266174 545134 305618
rect 544514 265938 544546 266174
rect 544782 265938 544866 266174
rect 545102 265938 545134 266174
rect 544514 265854 545134 265938
rect 544514 265618 544546 265854
rect 544782 265618 544866 265854
rect 545102 265618 545134 265854
rect 544514 226174 545134 265618
rect 544514 225938 544546 226174
rect 544782 225938 544866 226174
rect 545102 225938 545134 226174
rect 544514 225854 545134 225938
rect 544514 225618 544546 225854
rect 544782 225618 544866 225854
rect 545102 225618 545134 225854
rect 544514 186174 545134 225618
rect 544514 185938 544546 186174
rect 544782 185938 544866 186174
rect 545102 185938 545134 186174
rect 544514 185854 545134 185938
rect 544514 185618 544546 185854
rect 544782 185618 544866 185854
rect 545102 185618 545134 185854
rect 544514 146174 545134 185618
rect 544514 145938 544546 146174
rect 544782 145938 544866 146174
rect 545102 145938 545134 146174
rect 544514 145854 545134 145938
rect 544514 145618 544546 145854
rect 544782 145618 544866 145854
rect 545102 145618 545134 145854
rect 544514 106174 545134 145618
rect 544514 105938 544546 106174
rect 544782 105938 544866 106174
rect 545102 105938 545134 106174
rect 544514 105854 545134 105938
rect 544514 105618 544546 105854
rect 544782 105618 544866 105854
rect 545102 105618 545134 105854
rect 544514 66174 545134 105618
rect 544514 65938 544546 66174
rect 544782 65938 544866 66174
rect 545102 65938 545134 66174
rect 544514 65854 545134 65938
rect 544514 65618 544546 65854
rect 544782 65618 544866 65854
rect 545102 65618 545134 65854
rect 544514 26174 545134 65618
rect 544514 25938 544546 26174
rect 544782 25938 544866 26174
rect 545102 25938 545134 26174
rect 544514 25854 545134 25938
rect 544514 25618 544546 25854
rect 544782 25618 544866 25854
rect 545102 25618 545134 25854
rect 544514 -3226 545134 25618
rect 544514 -3462 544546 -3226
rect 544782 -3462 544866 -3226
rect 545102 -3462 545134 -3226
rect 544514 -3546 545134 -3462
rect 544514 -3782 544546 -3546
rect 544782 -3782 544866 -3546
rect 545102 -3782 545134 -3546
rect 544514 -3814 545134 -3782
rect 548234 669894 548854 709082
rect 548234 669658 548266 669894
rect 548502 669658 548586 669894
rect 548822 669658 548854 669894
rect 548234 669574 548854 669658
rect 548234 669338 548266 669574
rect 548502 669338 548586 669574
rect 548822 669338 548854 669574
rect 548234 629894 548854 669338
rect 548234 629658 548266 629894
rect 548502 629658 548586 629894
rect 548822 629658 548854 629894
rect 548234 629574 548854 629658
rect 548234 629338 548266 629574
rect 548502 629338 548586 629574
rect 548822 629338 548854 629574
rect 548234 589894 548854 629338
rect 548234 589658 548266 589894
rect 548502 589658 548586 589894
rect 548822 589658 548854 589894
rect 548234 589574 548854 589658
rect 548234 589338 548266 589574
rect 548502 589338 548586 589574
rect 548822 589338 548854 589574
rect 548234 549894 548854 589338
rect 548234 549658 548266 549894
rect 548502 549658 548586 549894
rect 548822 549658 548854 549894
rect 548234 549574 548854 549658
rect 548234 549338 548266 549574
rect 548502 549338 548586 549574
rect 548822 549338 548854 549574
rect 548234 509894 548854 549338
rect 548234 509658 548266 509894
rect 548502 509658 548586 509894
rect 548822 509658 548854 509894
rect 548234 509574 548854 509658
rect 548234 509338 548266 509574
rect 548502 509338 548586 509574
rect 548822 509338 548854 509574
rect 548234 469894 548854 509338
rect 548234 469658 548266 469894
rect 548502 469658 548586 469894
rect 548822 469658 548854 469894
rect 548234 469574 548854 469658
rect 548234 469338 548266 469574
rect 548502 469338 548586 469574
rect 548822 469338 548854 469574
rect 548234 429894 548854 469338
rect 548234 429658 548266 429894
rect 548502 429658 548586 429894
rect 548822 429658 548854 429894
rect 548234 429574 548854 429658
rect 548234 429338 548266 429574
rect 548502 429338 548586 429574
rect 548822 429338 548854 429574
rect 548234 389894 548854 429338
rect 548234 389658 548266 389894
rect 548502 389658 548586 389894
rect 548822 389658 548854 389894
rect 548234 389574 548854 389658
rect 548234 389338 548266 389574
rect 548502 389338 548586 389574
rect 548822 389338 548854 389574
rect 548234 349894 548854 389338
rect 548234 349658 548266 349894
rect 548502 349658 548586 349894
rect 548822 349658 548854 349894
rect 548234 349574 548854 349658
rect 548234 349338 548266 349574
rect 548502 349338 548586 349574
rect 548822 349338 548854 349574
rect 548234 309894 548854 349338
rect 548234 309658 548266 309894
rect 548502 309658 548586 309894
rect 548822 309658 548854 309894
rect 548234 309574 548854 309658
rect 548234 309338 548266 309574
rect 548502 309338 548586 309574
rect 548822 309338 548854 309574
rect 548234 269894 548854 309338
rect 548234 269658 548266 269894
rect 548502 269658 548586 269894
rect 548822 269658 548854 269894
rect 548234 269574 548854 269658
rect 548234 269338 548266 269574
rect 548502 269338 548586 269574
rect 548822 269338 548854 269574
rect 548234 229894 548854 269338
rect 548234 229658 548266 229894
rect 548502 229658 548586 229894
rect 548822 229658 548854 229894
rect 548234 229574 548854 229658
rect 548234 229338 548266 229574
rect 548502 229338 548586 229574
rect 548822 229338 548854 229574
rect 548234 189894 548854 229338
rect 548234 189658 548266 189894
rect 548502 189658 548586 189894
rect 548822 189658 548854 189894
rect 548234 189574 548854 189658
rect 548234 189338 548266 189574
rect 548502 189338 548586 189574
rect 548822 189338 548854 189574
rect 548234 149894 548854 189338
rect 548234 149658 548266 149894
rect 548502 149658 548586 149894
rect 548822 149658 548854 149894
rect 548234 149574 548854 149658
rect 548234 149338 548266 149574
rect 548502 149338 548586 149574
rect 548822 149338 548854 149574
rect 548234 109894 548854 149338
rect 548234 109658 548266 109894
rect 548502 109658 548586 109894
rect 548822 109658 548854 109894
rect 548234 109574 548854 109658
rect 548234 109338 548266 109574
rect 548502 109338 548586 109574
rect 548822 109338 548854 109574
rect 548234 69894 548854 109338
rect 548234 69658 548266 69894
rect 548502 69658 548586 69894
rect 548822 69658 548854 69894
rect 548234 69574 548854 69658
rect 548234 69338 548266 69574
rect 548502 69338 548586 69574
rect 548822 69338 548854 69574
rect 548234 29894 548854 69338
rect 548234 29658 548266 29894
rect 548502 29658 548586 29894
rect 548822 29658 548854 29894
rect 548234 29574 548854 29658
rect 548234 29338 548266 29574
rect 548502 29338 548586 29574
rect 548822 29338 548854 29574
rect 548234 -5146 548854 29338
rect 548234 -5382 548266 -5146
rect 548502 -5382 548586 -5146
rect 548822 -5382 548854 -5146
rect 548234 -5466 548854 -5382
rect 548234 -5702 548266 -5466
rect 548502 -5702 548586 -5466
rect 548822 -5702 548854 -5466
rect 548234 -5734 548854 -5702
rect 551954 673614 552574 711002
rect 571954 710598 572574 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 571954 710362 571986 710598
rect 572222 710362 572306 710598
rect 572542 710362 572574 710598
rect 571954 710278 572574 710362
rect 571954 710042 571986 710278
rect 572222 710042 572306 710278
rect 572542 710042 572574 710278
rect 568234 708678 568854 709670
rect 568234 708442 568266 708678
rect 568502 708442 568586 708678
rect 568822 708442 568854 708678
rect 568234 708358 568854 708442
rect 568234 708122 568266 708358
rect 568502 708122 568586 708358
rect 568822 708122 568854 708358
rect 564514 706758 565134 707750
rect 564514 706522 564546 706758
rect 564782 706522 564866 706758
rect 565102 706522 565134 706758
rect 564514 706438 565134 706522
rect 564514 706202 564546 706438
rect 564782 706202 564866 706438
rect 565102 706202 565134 706438
rect 551954 673378 551986 673614
rect 552222 673378 552306 673614
rect 552542 673378 552574 673614
rect 551954 673294 552574 673378
rect 551954 673058 551986 673294
rect 552222 673058 552306 673294
rect 552542 673058 552574 673294
rect 551954 633614 552574 673058
rect 551954 633378 551986 633614
rect 552222 633378 552306 633614
rect 552542 633378 552574 633614
rect 551954 633294 552574 633378
rect 551954 633058 551986 633294
rect 552222 633058 552306 633294
rect 552542 633058 552574 633294
rect 551954 593614 552574 633058
rect 551954 593378 551986 593614
rect 552222 593378 552306 593614
rect 552542 593378 552574 593614
rect 551954 593294 552574 593378
rect 551954 593058 551986 593294
rect 552222 593058 552306 593294
rect 552542 593058 552574 593294
rect 551954 553614 552574 593058
rect 551954 553378 551986 553614
rect 552222 553378 552306 553614
rect 552542 553378 552574 553614
rect 551954 553294 552574 553378
rect 551954 553058 551986 553294
rect 552222 553058 552306 553294
rect 552542 553058 552574 553294
rect 551954 513614 552574 553058
rect 551954 513378 551986 513614
rect 552222 513378 552306 513614
rect 552542 513378 552574 513614
rect 551954 513294 552574 513378
rect 551954 513058 551986 513294
rect 552222 513058 552306 513294
rect 552542 513058 552574 513294
rect 551954 473614 552574 513058
rect 551954 473378 551986 473614
rect 552222 473378 552306 473614
rect 552542 473378 552574 473614
rect 551954 473294 552574 473378
rect 551954 473058 551986 473294
rect 552222 473058 552306 473294
rect 552542 473058 552574 473294
rect 551954 433614 552574 473058
rect 551954 433378 551986 433614
rect 552222 433378 552306 433614
rect 552542 433378 552574 433614
rect 551954 433294 552574 433378
rect 551954 433058 551986 433294
rect 552222 433058 552306 433294
rect 552542 433058 552574 433294
rect 551954 393614 552574 433058
rect 551954 393378 551986 393614
rect 552222 393378 552306 393614
rect 552542 393378 552574 393614
rect 551954 393294 552574 393378
rect 551954 393058 551986 393294
rect 552222 393058 552306 393294
rect 552542 393058 552574 393294
rect 551954 353614 552574 393058
rect 551954 353378 551986 353614
rect 552222 353378 552306 353614
rect 552542 353378 552574 353614
rect 551954 353294 552574 353378
rect 551954 353058 551986 353294
rect 552222 353058 552306 353294
rect 552542 353058 552574 353294
rect 551954 313614 552574 353058
rect 551954 313378 551986 313614
rect 552222 313378 552306 313614
rect 552542 313378 552574 313614
rect 551954 313294 552574 313378
rect 551954 313058 551986 313294
rect 552222 313058 552306 313294
rect 552542 313058 552574 313294
rect 551954 273614 552574 313058
rect 551954 273378 551986 273614
rect 552222 273378 552306 273614
rect 552542 273378 552574 273614
rect 551954 273294 552574 273378
rect 551954 273058 551986 273294
rect 552222 273058 552306 273294
rect 552542 273058 552574 273294
rect 551954 233614 552574 273058
rect 551954 233378 551986 233614
rect 552222 233378 552306 233614
rect 552542 233378 552574 233614
rect 551954 233294 552574 233378
rect 551954 233058 551986 233294
rect 552222 233058 552306 233294
rect 552542 233058 552574 233294
rect 551954 193614 552574 233058
rect 551954 193378 551986 193614
rect 552222 193378 552306 193614
rect 552542 193378 552574 193614
rect 551954 193294 552574 193378
rect 551954 193058 551986 193294
rect 552222 193058 552306 193294
rect 552542 193058 552574 193294
rect 551954 153614 552574 193058
rect 551954 153378 551986 153614
rect 552222 153378 552306 153614
rect 552542 153378 552574 153614
rect 551954 153294 552574 153378
rect 551954 153058 551986 153294
rect 552222 153058 552306 153294
rect 552542 153058 552574 153294
rect 551954 113614 552574 153058
rect 551954 113378 551986 113614
rect 552222 113378 552306 113614
rect 552542 113378 552574 113614
rect 551954 113294 552574 113378
rect 551954 113058 551986 113294
rect 552222 113058 552306 113294
rect 552542 113058 552574 113294
rect 551954 73614 552574 113058
rect 551954 73378 551986 73614
rect 552222 73378 552306 73614
rect 552542 73378 552574 73614
rect 551954 73294 552574 73378
rect 551954 73058 551986 73294
rect 552222 73058 552306 73294
rect 552542 73058 552574 73294
rect 551954 33614 552574 73058
rect 551954 33378 551986 33614
rect 552222 33378 552306 33614
rect 552542 33378 552574 33614
rect 551954 33294 552574 33378
rect 551954 33058 551986 33294
rect 552222 33058 552306 33294
rect 552542 33058 552574 33294
rect 531954 -6342 531986 -6106
rect 532222 -6342 532306 -6106
rect 532542 -6342 532574 -6106
rect 531954 -6426 532574 -6342
rect 531954 -6662 531986 -6426
rect 532222 -6662 532306 -6426
rect 532542 -6662 532574 -6426
rect 531954 -7654 532574 -6662
rect 551954 -7066 552574 33058
rect 560794 704838 561414 705830
rect 560794 704602 560826 704838
rect 561062 704602 561146 704838
rect 561382 704602 561414 704838
rect 560794 704518 561414 704602
rect 560794 704282 560826 704518
rect 561062 704282 561146 704518
rect 561382 704282 561414 704518
rect 560794 682454 561414 704282
rect 560794 682218 560826 682454
rect 561062 682218 561146 682454
rect 561382 682218 561414 682454
rect 560794 682134 561414 682218
rect 560794 681898 560826 682134
rect 561062 681898 561146 682134
rect 561382 681898 561414 682134
rect 560794 642454 561414 681898
rect 560794 642218 560826 642454
rect 561062 642218 561146 642454
rect 561382 642218 561414 642454
rect 560794 642134 561414 642218
rect 560794 641898 560826 642134
rect 561062 641898 561146 642134
rect 561382 641898 561414 642134
rect 560794 602454 561414 641898
rect 560794 602218 560826 602454
rect 561062 602218 561146 602454
rect 561382 602218 561414 602454
rect 560794 602134 561414 602218
rect 560794 601898 560826 602134
rect 561062 601898 561146 602134
rect 561382 601898 561414 602134
rect 560794 562454 561414 601898
rect 560794 562218 560826 562454
rect 561062 562218 561146 562454
rect 561382 562218 561414 562454
rect 560794 562134 561414 562218
rect 560794 561898 560826 562134
rect 561062 561898 561146 562134
rect 561382 561898 561414 562134
rect 560794 522454 561414 561898
rect 560794 522218 560826 522454
rect 561062 522218 561146 522454
rect 561382 522218 561414 522454
rect 560794 522134 561414 522218
rect 560794 521898 560826 522134
rect 561062 521898 561146 522134
rect 561382 521898 561414 522134
rect 560794 482454 561414 521898
rect 560794 482218 560826 482454
rect 561062 482218 561146 482454
rect 561382 482218 561414 482454
rect 560794 482134 561414 482218
rect 560794 481898 560826 482134
rect 561062 481898 561146 482134
rect 561382 481898 561414 482134
rect 560794 442454 561414 481898
rect 560794 442218 560826 442454
rect 561062 442218 561146 442454
rect 561382 442218 561414 442454
rect 560794 442134 561414 442218
rect 560794 441898 560826 442134
rect 561062 441898 561146 442134
rect 561382 441898 561414 442134
rect 560794 402454 561414 441898
rect 560794 402218 560826 402454
rect 561062 402218 561146 402454
rect 561382 402218 561414 402454
rect 560794 402134 561414 402218
rect 560794 401898 560826 402134
rect 561062 401898 561146 402134
rect 561382 401898 561414 402134
rect 560794 362454 561414 401898
rect 560794 362218 560826 362454
rect 561062 362218 561146 362454
rect 561382 362218 561414 362454
rect 560794 362134 561414 362218
rect 560794 361898 560826 362134
rect 561062 361898 561146 362134
rect 561382 361898 561414 362134
rect 560794 322454 561414 361898
rect 560794 322218 560826 322454
rect 561062 322218 561146 322454
rect 561382 322218 561414 322454
rect 560794 322134 561414 322218
rect 560794 321898 560826 322134
rect 561062 321898 561146 322134
rect 561382 321898 561414 322134
rect 560794 282454 561414 321898
rect 560794 282218 560826 282454
rect 561062 282218 561146 282454
rect 561382 282218 561414 282454
rect 560794 282134 561414 282218
rect 560794 281898 560826 282134
rect 561062 281898 561146 282134
rect 561382 281898 561414 282134
rect 560794 242454 561414 281898
rect 560794 242218 560826 242454
rect 561062 242218 561146 242454
rect 561382 242218 561414 242454
rect 560794 242134 561414 242218
rect 560794 241898 560826 242134
rect 561062 241898 561146 242134
rect 561382 241898 561414 242134
rect 560794 202454 561414 241898
rect 560794 202218 560826 202454
rect 561062 202218 561146 202454
rect 561382 202218 561414 202454
rect 560794 202134 561414 202218
rect 560794 201898 560826 202134
rect 561062 201898 561146 202134
rect 561382 201898 561414 202134
rect 560794 162454 561414 201898
rect 560794 162218 560826 162454
rect 561062 162218 561146 162454
rect 561382 162218 561414 162454
rect 560794 162134 561414 162218
rect 560794 161898 560826 162134
rect 561062 161898 561146 162134
rect 561382 161898 561414 162134
rect 560794 122454 561414 161898
rect 560794 122218 560826 122454
rect 561062 122218 561146 122454
rect 561382 122218 561414 122454
rect 560794 122134 561414 122218
rect 560794 121898 560826 122134
rect 561062 121898 561146 122134
rect 561382 121898 561414 122134
rect 560794 82454 561414 121898
rect 560794 82218 560826 82454
rect 561062 82218 561146 82454
rect 561382 82218 561414 82454
rect 560794 82134 561414 82218
rect 560794 81898 560826 82134
rect 561062 81898 561146 82134
rect 561382 81898 561414 82134
rect 560794 42454 561414 81898
rect 560794 42218 560826 42454
rect 561062 42218 561146 42454
rect 561382 42218 561414 42454
rect 560794 42134 561414 42218
rect 560794 41898 560826 42134
rect 561062 41898 561146 42134
rect 561382 41898 561414 42134
rect 560794 2454 561414 41898
rect 560794 2218 560826 2454
rect 561062 2218 561146 2454
rect 561382 2218 561414 2454
rect 560794 2134 561414 2218
rect 560794 1898 560826 2134
rect 561062 1898 561146 2134
rect 561382 1898 561414 2134
rect 560794 -346 561414 1898
rect 560794 -582 560826 -346
rect 561062 -582 561146 -346
rect 561382 -582 561414 -346
rect 560794 -666 561414 -582
rect 560794 -902 560826 -666
rect 561062 -902 561146 -666
rect 561382 -902 561414 -666
rect 560794 -1894 561414 -902
rect 564514 686174 565134 706202
rect 564514 685938 564546 686174
rect 564782 685938 564866 686174
rect 565102 685938 565134 686174
rect 564514 685854 565134 685938
rect 564514 685618 564546 685854
rect 564782 685618 564866 685854
rect 565102 685618 565134 685854
rect 564514 646174 565134 685618
rect 564514 645938 564546 646174
rect 564782 645938 564866 646174
rect 565102 645938 565134 646174
rect 564514 645854 565134 645938
rect 564514 645618 564546 645854
rect 564782 645618 564866 645854
rect 565102 645618 565134 645854
rect 564514 606174 565134 645618
rect 564514 605938 564546 606174
rect 564782 605938 564866 606174
rect 565102 605938 565134 606174
rect 564514 605854 565134 605938
rect 564514 605618 564546 605854
rect 564782 605618 564866 605854
rect 565102 605618 565134 605854
rect 564514 566174 565134 605618
rect 564514 565938 564546 566174
rect 564782 565938 564866 566174
rect 565102 565938 565134 566174
rect 564514 565854 565134 565938
rect 564514 565618 564546 565854
rect 564782 565618 564866 565854
rect 565102 565618 565134 565854
rect 564514 526174 565134 565618
rect 564514 525938 564546 526174
rect 564782 525938 564866 526174
rect 565102 525938 565134 526174
rect 564514 525854 565134 525938
rect 564514 525618 564546 525854
rect 564782 525618 564866 525854
rect 565102 525618 565134 525854
rect 564514 486174 565134 525618
rect 564514 485938 564546 486174
rect 564782 485938 564866 486174
rect 565102 485938 565134 486174
rect 564514 485854 565134 485938
rect 564514 485618 564546 485854
rect 564782 485618 564866 485854
rect 565102 485618 565134 485854
rect 564514 446174 565134 485618
rect 564514 445938 564546 446174
rect 564782 445938 564866 446174
rect 565102 445938 565134 446174
rect 564514 445854 565134 445938
rect 564514 445618 564546 445854
rect 564782 445618 564866 445854
rect 565102 445618 565134 445854
rect 564514 406174 565134 445618
rect 564514 405938 564546 406174
rect 564782 405938 564866 406174
rect 565102 405938 565134 406174
rect 564514 405854 565134 405938
rect 564514 405618 564546 405854
rect 564782 405618 564866 405854
rect 565102 405618 565134 405854
rect 564514 366174 565134 405618
rect 564514 365938 564546 366174
rect 564782 365938 564866 366174
rect 565102 365938 565134 366174
rect 564514 365854 565134 365938
rect 564514 365618 564546 365854
rect 564782 365618 564866 365854
rect 565102 365618 565134 365854
rect 564514 326174 565134 365618
rect 564514 325938 564546 326174
rect 564782 325938 564866 326174
rect 565102 325938 565134 326174
rect 564514 325854 565134 325938
rect 564514 325618 564546 325854
rect 564782 325618 564866 325854
rect 565102 325618 565134 325854
rect 564514 286174 565134 325618
rect 564514 285938 564546 286174
rect 564782 285938 564866 286174
rect 565102 285938 565134 286174
rect 564514 285854 565134 285938
rect 564514 285618 564546 285854
rect 564782 285618 564866 285854
rect 565102 285618 565134 285854
rect 564514 246174 565134 285618
rect 564514 245938 564546 246174
rect 564782 245938 564866 246174
rect 565102 245938 565134 246174
rect 564514 245854 565134 245938
rect 564514 245618 564546 245854
rect 564782 245618 564866 245854
rect 565102 245618 565134 245854
rect 564514 206174 565134 245618
rect 564514 205938 564546 206174
rect 564782 205938 564866 206174
rect 565102 205938 565134 206174
rect 564514 205854 565134 205938
rect 564514 205618 564546 205854
rect 564782 205618 564866 205854
rect 565102 205618 565134 205854
rect 564514 166174 565134 205618
rect 564514 165938 564546 166174
rect 564782 165938 564866 166174
rect 565102 165938 565134 166174
rect 564514 165854 565134 165938
rect 564514 165618 564546 165854
rect 564782 165618 564866 165854
rect 565102 165618 565134 165854
rect 564514 126174 565134 165618
rect 564514 125938 564546 126174
rect 564782 125938 564866 126174
rect 565102 125938 565134 126174
rect 564514 125854 565134 125938
rect 564514 125618 564546 125854
rect 564782 125618 564866 125854
rect 565102 125618 565134 125854
rect 564514 86174 565134 125618
rect 564514 85938 564546 86174
rect 564782 85938 564866 86174
rect 565102 85938 565134 86174
rect 564514 85854 565134 85938
rect 564514 85618 564546 85854
rect 564782 85618 564866 85854
rect 565102 85618 565134 85854
rect 564514 46174 565134 85618
rect 564514 45938 564546 46174
rect 564782 45938 564866 46174
rect 565102 45938 565134 46174
rect 564514 45854 565134 45938
rect 564514 45618 564546 45854
rect 564782 45618 564866 45854
rect 565102 45618 565134 45854
rect 564514 6174 565134 45618
rect 564514 5938 564546 6174
rect 564782 5938 564866 6174
rect 565102 5938 565134 6174
rect 564514 5854 565134 5938
rect 564514 5618 564546 5854
rect 564782 5618 564866 5854
rect 565102 5618 565134 5854
rect 564514 -2266 565134 5618
rect 564514 -2502 564546 -2266
rect 564782 -2502 564866 -2266
rect 565102 -2502 565134 -2266
rect 564514 -2586 565134 -2502
rect 564514 -2822 564546 -2586
rect 564782 -2822 564866 -2586
rect 565102 -2822 565134 -2586
rect 564514 -3814 565134 -2822
rect 568234 689894 568854 708122
rect 568234 689658 568266 689894
rect 568502 689658 568586 689894
rect 568822 689658 568854 689894
rect 568234 689574 568854 689658
rect 568234 689338 568266 689574
rect 568502 689338 568586 689574
rect 568822 689338 568854 689574
rect 568234 649894 568854 689338
rect 568234 649658 568266 649894
rect 568502 649658 568586 649894
rect 568822 649658 568854 649894
rect 568234 649574 568854 649658
rect 568234 649338 568266 649574
rect 568502 649338 568586 649574
rect 568822 649338 568854 649574
rect 568234 609894 568854 649338
rect 568234 609658 568266 609894
rect 568502 609658 568586 609894
rect 568822 609658 568854 609894
rect 568234 609574 568854 609658
rect 568234 609338 568266 609574
rect 568502 609338 568586 609574
rect 568822 609338 568854 609574
rect 568234 569894 568854 609338
rect 568234 569658 568266 569894
rect 568502 569658 568586 569894
rect 568822 569658 568854 569894
rect 568234 569574 568854 569658
rect 568234 569338 568266 569574
rect 568502 569338 568586 569574
rect 568822 569338 568854 569574
rect 568234 529894 568854 569338
rect 568234 529658 568266 529894
rect 568502 529658 568586 529894
rect 568822 529658 568854 529894
rect 568234 529574 568854 529658
rect 568234 529338 568266 529574
rect 568502 529338 568586 529574
rect 568822 529338 568854 529574
rect 568234 489894 568854 529338
rect 568234 489658 568266 489894
rect 568502 489658 568586 489894
rect 568822 489658 568854 489894
rect 568234 489574 568854 489658
rect 568234 489338 568266 489574
rect 568502 489338 568586 489574
rect 568822 489338 568854 489574
rect 568234 449894 568854 489338
rect 568234 449658 568266 449894
rect 568502 449658 568586 449894
rect 568822 449658 568854 449894
rect 568234 449574 568854 449658
rect 568234 449338 568266 449574
rect 568502 449338 568586 449574
rect 568822 449338 568854 449574
rect 568234 409894 568854 449338
rect 568234 409658 568266 409894
rect 568502 409658 568586 409894
rect 568822 409658 568854 409894
rect 568234 409574 568854 409658
rect 568234 409338 568266 409574
rect 568502 409338 568586 409574
rect 568822 409338 568854 409574
rect 568234 369894 568854 409338
rect 568234 369658 568266 369894
rect 568502 369658 568586 369894
rect 568822 369658 568854 369894
rect 568234 369574 568854 369658
rect 568234 369338 568266 369574
rect 568502 369338 568586 369574
rect 568822 369338 568854 369574
rect 568234 329894 568854 369338
rect 568234 329658 568266 329894
rect 568502 329658 568586 329894
rect 568822 329658 568854 329894
rect 568234 329574 568854 329658
rect 568234 329338 568266 329574
rect 568502 329338 568586 329574
rect 568822 329338 568854 329574
rect 568234 289894 568854 329338
rect 568234 289658 568266 289894
rect 568502 289658 568586 289894
rect 568822 289658 568854 289894
rect 568234 289574 568854 289658
rect 568234 289338 568266 289574
rect 568502 289338 568586 289574
rect 568822 289338 568854 289574
rect 568234 249894 568854 289338
rect 568234 249658 568266 249894
rect 568502 249658 568586 249894
rect 568822 249658 568854 249894
rect 568234 249574 568854 249658
rect 568234 249338 568266 249574
rect 568502 249338 568586 249574
rect 568822 249338 568854 249574
rect 568234 209894 568854 249338
rect 568234 209658 568266 209894
rect 568502 209658 568586 209894
rect 568822 209658 568854 209894
rect 568234 209574 568854 209658
rect 568234 209338 568266 209574
rect 568502 209338 568586 209574
rect 568822 209338 568854 209574
rect 568234 169894 568854 209338
rect 568234 169658 568266 169894
rect 568502 169658 568586 169894
rect 568822 169658 568854 169894
rect 568234 169574 568854 169658
rect 568234 169338 568266 169574
rect 568502 169338 568586 169574
rect 568822 169338 568854 169574
rect 568234 129894 568854 169338
rect 568234 129658 568266 129894
rect 568502 129658 568586 129894
rect 568822 129658 568854 129894
rect 568234 129574 568854 129658
rect 568234 129338 568266 129574
rect 568502 129338 568586 129574
rect 568822 129338 568854 129574
rect 568234 89894 568854 129338
rect 568234 89658 568266 89894
rect 568502 89658 568586 89894
rect 568822 89658 568854 89894
rect 568234 89574 568854 89658
rect 568234 89338 568266 89574
rect 568502 89338 568586 89574
rect 568822 89338 568854 89574
rect 568234 49894 568854 89338
rect 568234 49658 568266 49894
rect 568502 49658 568586 49894
rect 568822 49658 568854 49894
rect 568234 49574 568854 49658
rect 568234 49338 568266 49574
rect 568502 49338 568586 49574
rect 568822 49338 568854 49574
rect 568234 9894 568854 49338
rect 568234 9658 568266 9894
rect 568502 9658 568586 9894
rect 568822 9658 568854 9894
rect 568234 9574 568854 9658
rect 568234 9338 568266 9574
rect 568502 9338 568586 9574
rect 568822 9338 568854 9574
rect 568234 -4186 568854 9338
rect 568234 -4422 568266 -4186
rect 568502 -4422 568586 -4186
rect 568822 -4422 568854 -4186
rect 568234 -4506 568854 -4422
rect 568234 -4742 568266 -4506
rect 568502 -4742 568586 -4506
rect 568822 -4742 568854 -4506
rect 568234 -5734 568854 -4742
rect 571954 693614 572574 710042
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 571954 693378 571986 693614
rect 572222 693378 572306 693614
rect 572542 693378 572574 693614
rect 571954 693294 572574 693378
rect 571954 693058 571986 693294
rect 572222 693058 572306 693294
rect 572542 693058 572574 693294
rect 571954 653614 572574 693058
rect 571954 653378 571986 653614
rect 572222 653378 572306 653614
rect 572542 653378 572574 653614
rect 571954 653294 572574 653378
rect 571954 653058 571986 653294
rect 572222 653058 572306 653294
rect 572542 653058 572574 653294
rect 571954 613614 572574 653058
rect 571954 613378 571986 613614
rect 572222 613378 572306 613614
rect 572542 613378 572574 613614
rect 571954 613294 572574 613378
rect 571954 613058 571986 613294
rect 572222 613058 572306 613294
rect 572542 613058 572574 613294
rect 571954 573614 572574 613058
rect 571954 573378 571986 573614
rect 572222 573378 572306 573614
rect 572542 573378 572574 573614
rect 571954 573294 572574 573378
rect 571954 573058 571986 573294
rect 572222 573058 572306 573294
rect 572542 573058 572574 573294
rect 571954 533614 572574 573058
rect 571954 533378 571986 533614
rect 572222 533378 572306 533614
rect 572542 533378 572574 533614
rect 571954 533294 572574 533378
rect 571954 533058 571986 533294
rect 572222 533058 572306 533294
rect 572542 533058 572574 533294
rect 571954 493614 572574 533058
rect 571954 493378 571986 493614
rect 572222 493378 572306 493614
rect 572542 493378 572574 493614
rect 571954 493294 572574 493378
rect 571954 493058 571986 493294
rect 572222 493058 572306 493294
rect 572542 493058 572574 493294
rect 571954 453614 572574 493058
rect 571954 453378 571986 453614
rect 572222 453378 572306 453614
rect 572542 453378 572574 453614
rect 571954 453294 572574 453378
rect 571954 453058 571986 453294
rect 572222 453058 572306 453294
rect 572542 453058 572574 453294
rect 571954 413614 572574 453058
rect 571954 413378 571986 413614
rect 572222 413378 572306 413614
rect 572542 413378 572574 413614
rect 571954 413294 572574 413378
rect 571954 413058 571986 413294
rect 572222 413058 572306 413294
rect 572542 413058 572574 413294
rect 571954 373614 572574 413058
rect 571954 373378 571986 373614
rect 572222 373378 572306 373614
rect 572542 373378 572574 373614
rect 571954 373294 572574 373378
rect 571954 373058 571986 373294
rect 572222 373058 572306 373294
rect 572542 373058 572574 373294
rect 571954 333614 572574 373058
rect 571954 333378 571986 333614
rect 572222 333378 572306 333614
rect 572542 333378 572574 333614
rect 571954 333294 572574 333378
rect 571954 333058 571986 333294
rect 572222 333058 572306 333294
rect 572542 333058 572574 333294
rect 571954 293614 572574 333058
rect 571954 293378 571986 293614
rect 572222 293378 572306 293614
rect 572542 293378 572574 293614
rect 571954 293294 572574 293378
rect 571954 293058 571986 293294
rect 572222 293058 572306 293294
rect 572542 293058 572574 293294
rect 571954 253614 572574 293058
rect 571954 253378 571986 253614
rect 572222 253378 572306 253614
rect 572542 253378 572574 253614
rect 571954 253294 572574 253378
rect 571954 253058 571986 253294
rect 572222 253058 572306 253294
rect 572542 253058 572574 253294
rect 571954 213614 572574 253058
rect 571954 213378 571986 213614
rect 572222 213378 572306 213614
rect 572542 213378 572574 213614
rect 571954 213294 572574 213378
rect 571954 213058 571986 213294
rect 572222 213058 572306 213294
rect 572542 213058 572574 213294
rect 571954 173614 572574 213058
rect 571954 173378 571986 173614
rect 572222 173378 572306 173614
rect 572542 173378 572574 173614
rect 571954 173294 572574 173378
rect 571954 173058 571986 173294
rect 572222 173058 572306 173294
rect 572542 173058 572574 173294
rect 571954 133614 572574 173058
rect 571954 133378 571986 133614
rect 572222 133378 572306 133614
rect 572542 133378 572574 133614
rect 571954 133294 572574 133378
rect 571954 133058 571986 133294
rect 572222 133058 572306 133294
rect 572542 133058 572574 133294
rect 571954 93614 572574 133058
rect 571954 93378 571986 93614
rect 572222 93378 572306 93614
rect 572542 93378 572574 93614
rect 571954 93294 572574 93378
rect 571954 93058 571986 93294
rect 572222 93058 572306 93294
rect 572542 93058 572574 93294
rect 571954 53614 572574 93058
rect 571954 53378 571986 53614
rect 572222 53378 572306 53614
rect 572542 53378 572574 53614
rect 571954 53294 572574 53378
rect 571954 53058 571986 53294
rect 572222 53058 572306 53294
rect 572542 53058 572574 53294
rect 571954 13614 572574 53058
rect 571954 13378 571986 13614
rect 572222 13378 572306 13614
rect 572542 13378 572574 13614
rect 571954 13294 572574 13378
rect 571954 13058 571986 13294
rect 572222 13058 572306 13294
rect 572542 13058 572574 13294
rect 551954 -7302 551986 -7066
rect 552222 -7302 552306 -7066
rect 552542 -7302 552574 -7066
rect 551954 -7386 552574 -7302
rect 551954 -7622 551986 -7386
rect 552222 -7622 552306 -7386
rect 552542 -7622 552574 -7386
rect 551954 -7654 552574 -7622
rect 571954 -6106 572574 13058
rect 580794 705798 581414 705830
rect 580794 705562 580826 705798
rect 581062 705562 581146 705798
rect 581382 705562 581414 705798
rect 580794 705478 581414 705562
rect 580794 705242 580826 705478
rect 581062 705242 581146 705478
rect 581382 705242 581414 705478
rect 580794 662454 581414 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 580794 662218 580826 662454
rect 581062 662218 581146 662454
rect 581382 662218 581414 662454
rect 580794 662134 581414 662218
rect 580794 661898 580826 662134
rect 581062 661898 581146 662134
rect 581382 661898 581414 662134
rect 580794 622454 581414 661898
rect 580794 622218 580826 622454
rect 581062 622218 581146 622454
rect 581382 622218 581414 622454
rect 580794 622134 581414 622218
rect 580794 621898 580826 622134
rect 581062 621898 581146 622134
rect 581382 621898 581414 622134
rect 580794 582454 581414 621898
rect 580794 582218 580826 582454
rect 581062 582218 581146 582454
rect 581382 582218 581414 582454
rect 580794 582134 581414 582218
rect 580794 581898 580826 582134
rect 581062 581898 581146 582134
rect 581382 581898 581414 582134
rect 580794 542454 581414 581898
rect 580794 542218 580826 542454
rect 581062 542218 581146 542454
rect 581382 542218 581414 542454
rect 580794 542134 581414 542218
rect 580794 541898 580826 542134
rect 581062 541898 581146 542134
rect 581382 541898 581414 542134
rect 580794 502454 581414 541898
rect 580794 502218 580826 502454
rect 581062 502218 581146 502454
rect 581382 502218 581414 502454
rect 580794 502134 581414 502218
rect 580794 501898 580826 502134
rect 581062 501898 581146 502134
rect 581382 501898 581414 502134
rect 580794 462454 581414 501898
rect 580794 462218 580826 462454
rect 581062 462218 581146 462454
rect 581382 462218 581414 462454
rect 580794 462134 581414 462218
rect 580794 461898 580826 462134
rect 581062 461898 581146 462134
rect 581382 461898 581414 462134
rect 580794 422454 581414 461898
rect 580794 422218 580826 422454
rect 581062 422218 581146 422454
rect 581382 422218 581414 422454
rect 580794 422134 581414 422218
rect 580794 421898 580826 422134
rect 581062 421898 581146 422134
rect 581382 421898 581414 422134
rect 580794 382454 581414 421898
rect 580794 382218 580826 382454
rect 581062 382218 581146 382454
rect 581382 382218 581414 382454
rect 580794 382134 581414 382218
rect 580794 381898 580826 382134
rect 581062 381898 581146 382134
rect 581382 381898 581414 382134
rect 580794 342454 581414 381898
rect 580794 342218 580826 342454
rect 581062 342218 581146 342454
rect 581382 342218 581414 342454
rect 580794 342134 581414 342218
rect 580794 341898 580826 342134
rect 581062 341898 581146 342134
rect 581382 341898 581414 342134
rect 580794 302454 581414 341898
rect 580794 302218 580826 302454
rect 581062 302218 581146 302454
rect 581382 302218 581414 302454
rect 580794 302134 581414 302218
rect 580794 301898 580826 302134
rect 581062 301898 581146 302134
rect 581382 301898 581414 302134
rect 580794 262454 581414 301898
rect 580794 262218 580826 262454
rect 581062 262218 581146 262454
rect 581382 262218 581414 262454
rect 580794 262134 581414 262218
rect 580794 261898 580826 262134
rect 581062 261898 581146 262134
rect 581382 261898 581414 262134
rect 580794 222454 581414 261898
rect 580794 222218 580826 222454
rect 581062 222218 581146 222454
rect 581382 222218 581414 222454
rect 580794 222134 581414 222218
rect 580794 221898 580826 222134
rect 581062 221898 581146 222134
rect 581382 221898 581414 222134
rect 580794 182454 581414 221898
rect 580794 182218 580826 182454
rect 581062 182218 581146 182454
rect 581382 182218 581414 182454
rect 580794 182134 581414 182218
rect 580794 181898 580826 182134
rect 581062 181898 581146 182134
rect 581382 181898 581414 182134
rect 580794 142454 581414 181898
rect 580794 142218 580826 142454
rect 581062 142218 581146 142454
rect 581382 142218 581414 142454
rect 580794 142134 581414 142218
rect 580794 141898 580826 142134
rect 581062 141898 581146 142134
rect 581382 141898 581414 142134
rect 580794 102454 581414 141898
rect 580794 102218 580826 102454
rect 581062 102218 581146 102454
rect 581382 102218 581414 102454
rect 580794 102134 581414 102218
rect 580794 101898 580826 102134
rect 581062 101898 581146 102134
rect 581382 101898 581414 102134
rect 580794 62454 581414 101898
rect 580794 62218 580826 62454
rect 581062 62218 581146 62454
rect 581382 62218 581414 62454
rect 580794 62134 581414 62218
rect 580794 61898 580826 62134
rect 581062 61898 581146 62134
rect 581382 61898 581414 62134
rect 580794 22454 581414 61898
rect 580794 22218 580826 22454
rect 581062 22218 581146 22454
rect 581382 22218 581414 22454
rect 580794 22134 581414 22218
rect 580794 21898 580826 22134
rect 581062 21898 581146 22134
rect 581382 21898 581414 22134
rect 580794 -1306 581414 21898
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 682454 585930 704282
rect 585310 682218 585342 682454
rect 585578 682218 585662 682454
rect 585898 682218 585930 682454
rect 585310 682134 585930 682218
rect 585310 681898 585342 682134
rect 585578 681898 585662 682134
rect 585898 681898 585930 682134
rect 585310 642454 585930 681898
rect 585310 642218 585342 642454
rect 585578 642218 585662 642454
rect 585898 642218 585930 642454
rect 585310 642134 585930 642218
rect 585310 641898 585342 642134
rect 585578 641898 585662 642134
rect 585898 641898 585930 642134
rect 585310 602454 585930 641898
rect 585310 602218 585342 602454
rect 585578 602218 585662 602454
rect 585898 602218 585930 602454
rect 585310 602134 585930 602218
rect 585310 601898 585342 602134
rect 585578 601898 585662 602134
rect 585898 601898 585930 602134
rect 585310 562454 585930 601898
rect 585310 562218 585342 562454
rect 585578 562218 585662 562454
rect 585898 562218 585930 562454
rect 585310 562134 585930 562218
rect 585310 561898 585342 562134
rect 585578 561898 585662 562134
rect 585898 561898 585930 562134
rect 585310 522454 585930 561898
rect 585310 522218 585342 522454
rect 585578 522218 585662 522454
rect 585898 522218 585930 522454
rect 585310 522134 585930 522218
rect 585310 521898 585342 522134
rect 585578 521898 585662 522134
rect 585898 521898 585930 522134
rect 585310 482454 585930 521898
rect 585310 482218 585342 482454
rect 585578 482218 585662 482454
rect 585898 482218 585930 482454
rect 585310 482134 585930 482218
rect 585310 481898 585342 482134
rect 585578 481898 585662 482134
rect 585898 481898 585930 482134
rect 585310 442454 585930 481898
rect 585310 442218 585342 442454
rect 585578 442218 585662 442454
rect 585898 442218 585930 442454
rect 585310 442134 585930 442218
rect 585310 441898 585342 442134
rect 585578 441898 585662 442134
rect 585898 441898 585930 442134
rect 585310 402454 585930 441898
rect 585310 402218 585342 402454
rect 585578 402218 585662 402454
rect 585898 402218 585930 402454
rect 585310 402134 585930 402218
rect 585310 401898 585342 402134
rect 585578 401898 585662 402134
rect 585898 401898 585930 402134
rect 585310 362454 585930 401898
rect 585310 362218 585342 362454
rect 585578 362218 585662 362454
rect 585898 362218 585930 362454
rect 585310 362134 585930 362218
rect 585310 361898 585342 362134
rect 585578 361898 585662 362134
rect 585898 361898 585930 362134
rect 585310 322454 585930 361898
rect 585310 322218 585342 322454
rect 585578 322218 585662 322454
rect 585898 322218 585930 322454
rect 585310 322134 585930 322218
rect 585310 321898 585342 322134
rect 585578 321898 585662 322134
rect 585898 321898 585930 322134
rect 585310 282454 585930 321898
rect 585310 282218 585342 282454
rect 585578 282218 585662 282454
rect 585898 282218 585930 282454
rect 585310 282134 585930 282218
rect 585310 281898 585342 282134
rect 585578 281898 585662 282134
rect 585898 281898 585930 282134
rect 585310 242454 585930 281898
rect 585310 242218 585342 242454
rect 585578 242218 585662 242454
rect 585898 242218 585930 242454
rect 585310 242134 585930 242218
rect 585310 241898 585342 242134
rect 585578 241898 585662 242134
rect 585898 241898 585930 242134
rect 585310 202454 585930 241898
rect 585310 202218 585342 202454
rect 585578 202218 585662 202454
rect 585898 202218 585930 202454
rect 585310 202134 585930 202218
rect 585310 201898 585342 202134
rect 585578 201898 585662 202134
rect 585898 201898 585930 202134
rect 585310 162454 585930 201898
rect 585310 162218 585342 162454
rect 585578 162218 585662 162454
rect 585898 162218 585930 162454
rect 585310 162134 585930 162218
rect 585310 161898 585342 162134
rect 585578 161898 585662 162134
rect 585898 161898 585930 162134
rect 585310 122454 585930 161898
rect 585310 122218 585342 122454
rect 585578 122218 585662 122454
rect 585898 122218 585930 122454
rect 585310 122134 585930 122218
rect 585310 121898 585342 122134
rect 585578 121898 585662 122134
rect 585898 121898 585930 122134
rect 585310 82454 585930 121898
rect 585310 82218 585342 82454
rect 585578 82218 585662 82454
rect 585898 82218 585930 82454
rect 585310 82134 585930 82218
rect 585310 81898 585342 82134
rect 585578 81898 585662 82134
rect 585898 81898 585930 82134
rect 585310 42454 585930 81898
rect 585310 42218 585342 42454
rect 585578 42218 585662 42454
rect 585898 42218 585930 42454
rect 585310 42134 585930 42218
rect 585310 41898 585342 42134
rect 585578 41898 585662 42134
rect 585898 41898 585930 42134
rect 585310 2454 585930 41898
rect 585310 2218 585342 2454
rect 585578 2218 585662 2454
rect 585898 2218 585930 2454
rect 585310 2134 585930 2218
rect 585310 1898 585342 2134
rect 585578 1898 585662 2134
rect 585898 1898 585930 2134
rect 585310 -346 585930 1898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 662454 586890 705242
rect 586270 662218 586302 662454
rect 586538 662218 586622 662454
rect 586858 662218 586890 662454
rect 586270 662134 586890 662218
rect 586270 661898 586302 662134
rect 586538 661898 586622 662134
rect 586858 661898 586890 662134
rect 586270 622454 586890 661898
rect 586270 622218 586302 622454
rect 586538 622218 586622 622454
rect 586858 622218 586890 622454
rect 586270 622134 586890 622218
rect 586270 621898 586302 622134
rect 586538 621898 586622 622134
rect 586858 621898 586890 622134
rect 586270 582454 586890 621898
rect 586270 582218 586302 582454
rect 586538 582218 586622 582454
rect 586858 582218 586890 582454
rect 586270 582134 586890 582218
rect 586270 581898 586302 582134
rect 586538 581898 586622 582134
rect 586858 581898 586890 582134
rect 586270 542454 586890 581898
rect 586270 542218 586302 542454
rect 586538 542218 586622 542454
rect 586858 542218 586890 542454
rect 586270 542134 586890 542218
rect 586270 541898 586302 542134
rect 586538 541898 586622 542134
rect 586858 541898 586890 542134
rect 586270 502454 586890 541898
rect 586270 502218 586302 502454
rect 586538 502218 586622 502454
rect 586858 502218 586890 502454
rect 586270 502134 586890 502218
rect 586270 501898 586302 502134
rect 586538 501898 586622 502134
rect 586858 501898 586890 502134
rect 586270 462454 586890 501898
rect 586270 462218 586302 462454
rect 586538 462218 586622 462454
rect 586858 462218 586890 462454
rect 586270 462134 586890 462218
rect 586270 461898 586302 462134
rect 586538 461898 586622 462134
rect 586858 461898 586890 462134
rect 586270 422454 586890 461898
rect 586270 422218 586302 422454
rect 586538 422218 586622 422454
rect 586858 422218 586890 422454
rect 586270 422134 586890 422218
rect 586270 421898 586302 422134
rect 586538 421898 586622 422134
rect 586858 421898 586890 422134
rect 586270 382454 586890 421898
rect 586270 382218 586302 382454
rect 586538 382218 586622 382454
rect 586858 382218 586890 382454
rect 586270 382134 586890 382218
rect 586270 381898 586302 382134
rect 586538 381898 586622 382134
rect 586858 381898 586890 382134
rect 586270 342454 586890 381898
rect 586270 342218 586302 342454
rect 586538 342218 586622 342454
rect 586858 342218 586890 342454
rect 586270 342134 586890 342218
rect 586270 341898 586302 342134
rect 586538 341898 586622 342134
rect 586858 341898 586890 342134
rect 586270 302454 586890 341898
rect 586270 302218 586302 302454
rect 586538 302218 586622 302454
rect 586858 302218 586890 302454
rect 586270 302134 586890 302218
rect 586270 301898 586302 302134
rect 586538 301898 586622 302134
rect 586858 301898 586890 302134
rect 586270 262454 586890 301898
rect 586270 262218 586302 262454
rect 586538 262218 586622 262454
rect 586858 262218 586890 262454
rect 586270 262134 586890 262218
rect 586270 261898 586302 262134
rect 586538 261898 586622 262134
rect 586858 261898 586890 262134
rect 586270 222454 586890 261898
rect 586270 222218 586302 222454
rect 586538 222218 586622 222454
rect 586858 222218 586890 222454
rect 586270 222134 586890 222218
rect 586270 221898 586302 222134
rect 586538 221898 586622 222134
rect 586858 221898 586890 222134
rect 586270 182454 586890 221898
rect 586270 182218 586302 182454
rect 586538 182218 586622 182454
rect 586858 182218 586890 182454
rect 586270 182134 586890 182218
rect 586270 181898 586302 182134
rect 586538 181898 586622 182134
rect 586858 181898 586890 182134
rect 586270 142454 586890 181898
rect 586270 142218 586302 142454
rect 586538 142218 586622 142454
rect 586858 142218 586890 142454
rect 586270 142134 586890 142218
rect 586270 141898 586302 142134
rect 586538 141898 586622 142134
rect 586858 141898 586890 142134
rect 586270 102454 586890 141898
rect 586270 102218 586302 102454
rect 586538 102218 586622 102454
rect 586858 102218 586890 102454
rect 586270 102134 586890 102218
rect 586270 101898 586302 102134
rect 586538 101898 586622 102134
rect 586858 101898 586890 102134
rect 586270 62454 586890 101898
rect 586270 62218 586302 62454
rect 586538 62218 586622 62454
rect 586858 62218 586890 62454
rect 586270 62134 586890 62218
rect 586270 61898 586302 62134
rect 586538 61898 586622 62134
rect 586858 61898 586890 62134
rect 586270 22454 586890 61898
rect 586270 22218 586302 22454
rect 586538 22218 586622 22454
rect 586858 22218 586890 22454
rect 586270 22134 586890 22218
rect 586270 21898 586302 22134
rect 586538 21898 586622 22134
rect 586858 21898 586890 22134
rect 580794 -1542 580826 -1306
rect 581062 -1542 581146 -1306
rect 581382 -1542 581414 -1306
rect 580794 -1626 581414 -1542
rect 580794 -1862 580826 -1626
rect 581062 -1862 581146 -1626
rect 581382 -1862 581414 -1626
rect 580794 -1894 581414 -1862
rect 586270 -1306 586890 21898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 686174 587850 706202
rect 587230 685938 587262 686174
rect 587498 685938 587582 686174
rect 587818 685938 587850 686174
rect 587230 685854 587850 685938
rect 587230 685618 587262 685854
rect 587498 685618 587582 685854
rect 587818 685618 587850 685854
rect 587230 646174 587850 685618
rect 587230 645938 587262 646174
rect 587498 645938 587582 646174
rect 587818 645938 587850 646174
rect 587230 645854 587850 645938
rect 587230 645618 587262 645854
rect 587498 645618 587582 645854
rect 587818 645618 587850 645854
rect 587230 606174 587850 645618
rect 587230 605938 587262 606174
rect 587498 605938 587582 606174
rect 587818 605938 587850 606174
rect 587230 605854 587850 605938
rect 587230 605618 587262 605854
rect 587498 605618 587582 605854
rect 587818 605618 587850 605854
rect 587230 566174 587850 605618
rect 587230 565938 587262 566174
rect 587498 565938 587582 566174
rect 587818 565938 587850 566174
rect 587230 565854 587850 565938
rect 587230 565618 587262 565854
rect 587498 565618 587582 565854
rect 587818 565618 587850 565854
rect 587230 526174 587850 565618
rect 587230 525938 587262 526174
rect 587498 525938 587582 526174
rect 587818 525938 587850 526174
rect 587230 525854 587850 525938
rect 587230 525618 587262 525854
rect 587498 525618 587582 525854
rect 587818 525618 587850 525854
rect 587230 486174 587850 525618
rect 587230 485938 587262 486174
rect 587498 485938 587582 486174
rect 587818 485938 587850 486174
rect 587230 485854 587850 485938
rect 587230 485618 587262 485854
rect 587498 485618 587582 485854
rect 587818 485618 587850 485854
rect 587230 446174 587850 485618
rect 587230 445938 587262 446174
rect 587498 445938 587582 446174
rect 587818 445938 587850 446174
rect 587230 445854 587850 445938
rect 587230 445618 587262 445854
rect 587498 445618 587582 445854
rect 587818 445618 587850 445854
rect 587230 406174 587850 445618
rect 587230 405938 587262 406174
rect 587498 405938 587582 406174
rect 587818 405938 587850 406174
rect 587230 405854 587850 405938
rect 587230 405618 587262 405854
rect 587498 405618 587582 405854
rect 587818 405618 587850 405854
rect 587230 366174 587850 405618
rect 587230 365938 587262 366174
rect 587498 365938 587582 366174
rect 587818 365938 587850 366174
rect 587230 365854 587850 365938
rect 587230 365618 587262 365854
rect 587498 365618 587582 365854
rect 587818 365618 587850 365854
rect 587230 326174 587850 365618
rect 587230 325938 587262 326174
rect 587498 325938 587582 326174
rect 587818 325938 587850 326174
rect 587230 325854 587850 325938
rect 587230 325618 587262 325854
rect 587498 325618 587582 325854
rect 587818 325618 587850 325854
rect 587230 286174 587850 325618
rect 587230 285938 587262 286174
rect 587498 285938 587582 286174
rect 587818 285938 587850 286174
rect 587230 285854 587850 285938
rect 587230 285618 587262 285854
rect 587498 285618 587582 285854
rect 587818 285618 587850 285854
rect 587230 246174 587850 285618
rect 587230 245938 587262 246174
rect 587498 245938 587582 246174
rect 587818 245938 587850 246174
rect 587230 245854 587850 245938
rect 587230 245618 587262 245854
rect 587498 245618 587582 245854
rect 587818 245618 587850 245854
rect 587230 206174 587850 245618
rect 587230 205938 587262 206174
rect 587498 205938 587582 206174
rect 587818 205938 587850 206174
rect 587230 205854 587850 205938
rect 587230 205618 587262 205854
rect 587498 205618 587582 205854
rect 587818 205618 587850 205854
rect 587230 166174 587850 205618
rect 587230 165938 587262 166174
rect 587498 165938 587582 166174
rect 587818 165938 587850 166174
rect 587230 165854 587850 165938
rect 587230 165618 587262 165854
rect 587498 165618 587582 165854
rect 587818 165618 587850 165854
rect 587230 126174 587850 165618
rect 587230 125938 587262 126174
rect 587498 125938 587582 126174
rect 587818 125938 587850 126174
rect 587230 125854 587850 125938
rect 587230 125618 587262 125854
rect 587498 125618 587582 125854
rect 587818 125618 587850 125854
rect 587230 86174 587850 125618
rect 587230 85938 587262 86174
rect 587498 85938 587582 86174
rect 587818 85938 587850 86174
rect 587230 85854 587850 85938
rect 587230 85618 587262 85854
rect 587498 85618 587582 85854
rect 587818 85618 587850 85854
rect 587230 46174 587850 85618
rect 587230 45938 587262 46174
rect 587498 45938 587582 46174
rect 587818 45938 587850 46174
rect 587230 45854 587850 45938
rect 587230 45618 587262 45854
rect 587498 45618 587582 45854
rect 587818 45618 587850 45854
rect 587230 6174 587850 45618
rect 587230 5938 587262 6174
rect 587498 5938 587582 6174
rect 587818 5938 587850 6174
rect 587230 5854 587850 5938
rect 587230 5618 587262 5854
rect 587498 5618 587582 5854
rect 587818 5618 587850 5854
rect 587230 -2266 587850 5618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 666174 588810 707162
rect 588190 665938 588222 666174
rect 588458 665938 588542 666174
rect 588778 665938 588810 666174
rect 588190 665854 588810 665938
rect 588190 665618 588222 665854
rect 588458 665618 588542 665854
rect 588778 665618 588810 665854
rect 588190 626174 588810 665618
rect 588190 625938 588222 626174
rect 588458 625938 588542 626174
rect 588778 625938 588810 626174
rect 588190 625854 588810 625938
rect 588190 625618 588222 625854
rect 588458 625618 588542 625854
rect 588778 625618 588810 625854
rect 588190 586174 588810 625618
rect 588190 585938 588222 586174
rect 588458 585938 588542 586174
rect 588778 585938 588810 586174
rect 588190 585854 588810 585938
rect 588190 585618 588222 585854
rect 588458 585618 588542 585854
rect 588778 585618 588810 585854
rect 588190 546174 588810 585618
rect 588190 545938 588222 546174
rect 588458 545938 588542 546174
rect 588778 545938 588810 546174
rect 588190 545854 588810 545938
rect 588190 545618 588222 545854
rect 588458 545618 588542 545854
rect 588778 545618 588810 545854
rect 588190 506174 588810 545618
rect 588190 505938 588222 506174
rect 588458 505938 588542 506174
rect 588778 505938 588810 506174
rect 588190 505854 588810 505938
rect 588190 505618 588222 505854
rect 588458 505618 588542 505854
rect 588778 505618 588810 505854
rect 588190 466174 588810 505618
rect 588190 465938 588222 466174
rect 588458 465938 588542 466174
rect 588778 465938 588810 466174
rect 588190 465854 588810 465938
rect 588190 465618 588222 465854
rect 588458 465618 588542 465854
rect 588778 465618 588810 465854
rect 588190 426174 588810 465618
rect 588190 425938 588222 426174
rect 588458 425938 588542 426174
rect 588778 425938 588810 426174
rect 588190 425854 588810 425938
rect 588190 425618 588222 425854
rect 588458 425618 588542 425854
rect 588778 425618 588810 425854
rect 588190 386174 588810 425618
rect 588190 385938 588222 386174
rect 588458 385938 588542 386174
rect 588778 385938 588810 386174
rect 588190 385854 588810 385938
rect 588190 385618 588222 385854
rect 588458 385618 588542 385854
rect 588778 385618 588810 385854
rect 588190 346174 588810 385618
rect 588190 345938 588222 346174
rect 588458 345938 588542 346174
rect 588778 345938 588810 346174
rect 588190 345854 588810 345938
rect 588190 345618 588222 345854
rect 588458 345618 588542 345854
rect 588778 345618 588810 345854
rect 588190 306174 588810 345618
rect 588190 305938 588222 306174
rect 588458 305938 588542 306174
rect 588778 305938 588810 306174
rect 588190 305854 588810 305938
rect 588190 305618 588222 305854
rect 588458 305618 588542 305854
rect 588778 305618 588810 305854
rect 588190 266174 588810 305618
rect 588190 265938 588222 266174
rect 588458 265938 588542 266174
rect 588778 265938 588810 266174
rect 588190 265854 588810 265938
rect 588190 265618 588222 265854
rect 588458 265618 588542 265854
rect 588778 265618 588810 265854
rect 588190 226174 588810 265618
rect 588190 225938 588222 226174
rect 588458 225938 588542 226174
rect 588778 225938 588810 226174
rect 588190 225854 588810 225938
rect 588190 225618 588222 225854
rect 588458 225618 588542 225854
rect 588778 225618 588810 225854
rect 588190 186174 588810 225618
rect 588190 185938 588222 186174
rect 588458 185938 588542 186174
rect 588778 185938 588810 186174
rect 588190 185854 588810 185938
rect 588190 185618 588222 185854
rect 588458 185618 588542 185854
rect 588778 185618 588810 185854
rect 588190 146174 588810 185618
rect 588190 145938 588222 146174
rect 588458 145938 588542 146174
rect 588778 145938 588810 146174
rect 588190 145854 588810 145938
rect 588190 145618 588222 145854
rect 588458 145618 588542 145854
rect 588778 145618 588810 145854
rect 588190 106174 588810 145618
rect 588190 105938 588222 106174
rect 588458 105938 588542 106174
rect 588778 105938 588810 106174
rect 588190 105854 588810 105938
rect 588190 105618 588222 105854
rect 588458 105618 588542 105854
rect 588778 105618 588810 105854
rect 588190 66174 588810 105618
rect 588190 65938 588222 66174
rect 588458 65938 588542 66174
rect 588778 65938 588810 66174
rect 588190 65854 588810 65938
rect 588190 65618 588222 65854
rect 588458 65618 588542 65854
rect 588778 65618 588810 65854
rect 588190 26174 588810 65618
rect 588190 25938 588222 26174
rect 588458 25938 588542 26174
rect 588778 25938 588810 26174
rect 588190 25854 588810 25938
rect 588190 25618 588222 25854
rect 588458 25618 588542 25854
rect 588778 25618 588810 25854
rect 588190 -3226 588810 25618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 689894 589770 708122
rect 589150 689658 589182 689894
rect 589418 689658 589502 689894
rect 589738 689658 589770 689894
rect 589150 689574 589770 689658
rect 589150 689338 589182 689574
rect 589418 689338 589502 689574
rect 589738 689338 589770 689574
rect 589150 649894 589770 689338
rect 589150 649658 589182 649894
rect 589418 649658 589502 649894
rect 589738 649658 589770 649894
rect 589150 649574 589770 649658
rect 589150 649338 589182 649574
rect 589418 649338 589502 649574
rect 589738 649338 589770 649574
rect 589150 609894 589770 649338
rect 589150 609658 589182 609894
rect 589418 609658 589502 609894
rect 589738 609658 589770 609894
rect 589150 609574 589770 609658
rect 589150 609338 589182 609574
rect 589418 609338 589502 609574
rect 589738 609338 589770 609574
rect 589150 569894 589770 609338
rect 589150 569658 589182 569894
rect 589418 569658 589502 569894
rect 589738 569658 589770 569894
rect 589150 569574 589770 569658
rect 589150 569338 589182 569574
rect 589418 569338 589502 569574
rect 589738 569338 589770 569574
rect 589150 529894 589770 569338
rect 589150 529658 589182 529894
rect 589418 529658 589502 529894
rect 589738 529658 589770 529894
rect 589150 529574 589770 529658
rect 589150 529338 589182 529574
rect 589418 529338 589502 529574
rect 589738 529338 589770 529574
rect 589150 489894 589770 529338
rect 589150 489658 589182 489894
rect 589418 489658 589502 489894
rect 589738 489658 589770 489894
rect 589150 489574 589770 489658
rect 589150 489338 589182 489574
rect 589418 489338 589502 489574
rect 589738 489338 589770 489574
rect 589150 449894 589770 489338
rect 589150 449658 589182 449894
rect 589418 449658 589502 449894
rect 589738 449658 589770 449894
rect 589150 449574 589770 449658
rect 589150 449338 589182 449574
rect 589418 449338 589502 449574
rect 589738 449338 589770 449574
rect 589150 409894 589770 449338
rect 589150 409658 589182 409894
rect 589418 409658 589502 409894
rect 589738 409658 589770 409894
rect 589150 409574 589770 409658
rect 589150 409338 589182 409574
rect 589418 409338 589502 409574
rect 589738 409338 589770 409574
rect 589150 369894 589770 409338
rect 589150 369658 589182 369894
rect 589418 369658 589502 369894
rect 589738 369658 589770 369894
rect 589150 369574 589770 369658
rect 589150 369338 589182 369574
rect 589418 369338 589502 369574
rect 589738 369338 589770 369574
rect 589150 329894 589770 369338
rect 589150 329658 589182 329894
rect 589418 329658 589502 329894
rect 589738 329658 589770 329894
rect 589150 329574 589770 329658
rect 589150 329338 589182 329574
rect 589418 329338 589502 329574
rect 589738 329338 589770 329574
rect 589150 289894 589770 329338
rect 589150 289658 589182 289894
rect 589418 289658 589502 289894
rect 589738 289658 589770 289894
rect 589150 289574 589770 289658
rect 589150 289338 589182 289574
rect 589418 289338 589502 289574
rect 589738 289338 589770 289574
rect 589150 249894 589770 289338
rect 589150 249658 589182 249894
rect 589418 249658 589502 249894
rect 589738 249658 589770 249894
rect 589150 249574 589770 249658
rect 589150 249338 589182 249574
rect 589418 249338 589502 249574
rect 589738 249338 589770 249574
rect 589150 209894 589770 249338
rect 589150 209658 589182 209894
rect 589418 209658 589502 209894
rect 589738 209658 589770 209894
rect 589150 209574 589770 209658
rect 589150 209338 589182 209574
rect 589418 209338 589502 209574
rect 589738 209338 589770 209574
rect 589150 169894 589770 209338
rect 589150 169658 589182 169894
rect 589418 169658 589502 169894
rect 589738 169658 589770 169894
rect 589150 169574 589770 169658
rect 589150 169338 589182 169574
rect 589418 169338 589502 169574
rect 589738 169338 589770 169574
rect 589150 129894 589770 169338
rect 589150 129658 589182 129894
rect 589418 129658 589502 129894
rect 589738 129658 589770 129894
rect 589150 129574 589770 129658
rect 589150 129338 589182 129574
rect 589418 129338 589502 129574
rect 589738 129338 589770 129574
rect 589150 89894 589770 129338
rect 589150 89658 589182 89894
rect 589418 89658 589502 89894
rect 589738 89658 589770 89894
rect 589150 89574 589770 89658
rect 589150 89338 589182 89574
rect 589418 89338 589502 89574
rect 589738 89338 589770 89574
rect 589150 49894 589770 89338
rect 589150 49658 589182 49894
rect 589418 49658 589502 49894
rect 589738 49658 589770 49894
rect 589150 49574 589770 49658
rect 589150 49338 589182 49574
rect 589418 49338 589502 49574
rect 589738 49338 589770 49574
rect 589150 9894 589770 49338
rect 589150 9658 589182 9894
rect 589418 9658 589502 9894
rect 589738 9658 589770 9894
rect 589150 9574 589770 9658
rect 589150 9338 589182 9574
rect 589418 9338 589502 9574
rect 589738 9338 589770 9574
rect 589150 -4186 589770 9338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 669894 590730 709082
rect 590110 669658 590142 669894
rect 590378 669658 590462 669894
rect 590698 669658 590730 669894
rect 590110 669574 590730 669658
rect 590110 669338 590142 669574
rect 590378 669338 590462 669574
rect 590698 669338 590730 669574
rect 590110 629894 590730 669338
rect 590110 629658 590142 629894
rect 590378 629658 590462 629894
rect 590698 629658 590730 629894
rect 590110 629574 590730 629658
rect 590110 629338 590142 629574
rect 590378 629338 590462 629574
rect 590698 629338 590730 629574
rect 590110 589894 590730 629338
rect 590110 589658 590142 589894
rect 590378 589658 590462 589894
rect 590698 589658 590730 589894
rect 590110 589574 590730 589658
rect 590110 589338 590142 589574
rect 590378 589338 590462 589574
rect 590698 589338 590730 589574
rect 590110 549894 590730 589338
rect 590110 549658 590142 549894
rect 590378 549658 590462 549894
rect 590698 549658 590730 549894
rect 590110 549574 590730 549658
rect 590110 549338 590142 549574
rect 590378 549338 590462 549574
rect 590698 549338 590730 549574
rect 590110 509894 590730 549338
rect 590110 509658 590142 509894
rect 590378 509658 590462 509894
rect 590698 509658 590730 509894
rect 590110 509574 590730 509658
rect 590110 509338 590142 509574
rect 590378 509338 590462 509574
rect 590698 509338 590730 509574
rect 590110 469894 590730 509338
rect 590110 469658 590142 469894
rect 590378 469658 590462 469894
rect 590698 469658 590730 469894
rect 590110 469574 590730 469658
rect 590110 469338 590142 469574
rect 590378 469338 590462 469574
rect 590698 469338 590730 469574
rect 590110 429894 590730 469338
rect 590110 429658 590142 429894
rect 590378 429658 590462 429894
rect 590698 429658 590730 429894
rect 590110 429574 590730 429658
rect 590110 429338 590142 429574
rect 590378 429338 590462 429574
rect 590698 429338 590730 429574
rect 590110 389894 590730 429338
rect 590110 389658 590142 389894
rect 590378 389658 590462 389894
rect 590698 389658 590730 389894
rect 590110 389574 590730 389658
rect 590110 389338 590142 389574
rect 590378 389338 590462 389574
rect 590698 389338 590730 389574
rect 590110 349894 590730 389338
rect 590110 349658 590142 349894
rect 590378 349658 590462 349894
rect 590698 349658 590730 349894
rect 590110 349574 590730 349658
rect 590110 349338 590142 349574
rect 590378 349338 590462 349574
rect 590698 349338 590730 349574
rect 590110 309894 590730 349338
rect 590110 309658 590142 309894
rect 590378 309658 590462 309894
rect 590698 309658 590730 309894
rect 590110 309574 590730 309658
rect 590110 309338 590142 309574
rect 590378 309338 590462 309574
rect 590698 309338 590730 309574
rect 590110 269894 590730 309338
rect 590110 269658 590142 269894
rect 590378 269658 590462 269894
rect 590698 269658 590730 269894
rect 590110 269574 590730 269658
rect 590110 269338 590142 269574
rect 590378 269338 590462 269574
rect 590698 269338 590730 269574
rect 590110 229894 590730 269338
rect 590110 229658 590142 229894
rect 590378 229658 590462 229894
rect 590698 229658 590730 229894
rect 590110 229574 590730 229658
rect 590110 229338 590142 229574
rect 590378 229338 590462 229574
rect 590698 229338 590730 229574
rect 590110 189894 590730 229338
rect 590110 189658 590142 189894
rect 590378 189658 590462 189894
rect 590698 189658 590730 189894
rect 590110 189574 590730 189658
rect 590110 189338 590142 189574
rect 590378 189338 590462 189574
rect 590698 189338 590730 189574
rect 590110 149894 590730 189338
rect 590110 149658 590142 149894
rect 590378 149658 590462 149894
rect 590698 149658 590730 149894
rect 590110 149574 590730 149658
rect 590110 149338 590142 149574
rect 590378 149338 590462 149574
rect 590698 149338 590730 149574
rect 590110 109894 590730 149338
rect 590110 109658 590142 109894
rect 590378 109658 590462 109894
rect 590698 109658 590730 109894
rect 590110 109574 590730 109658
rect 590110 109338 590142 109574
rect 590378 109338 590462 109574
rect 590698 109338 590730 109574
rect 590110 69894 590730 109338
rect 590110 69658 590142 69894
rect 590378 69658 590462 69894
rect 590698 69658 590730 69894
rect 590110 69574 590730 69658
rect 590110 69338 590142 69574
rect 590378 69338 590462 69574
rect 590698 69338 590730 69574
rect 590110 29894 590730 69338
rect 590110 29658 590142 29894
rect 590378 29658 590462 29894
rect 590698 29658 590730 29894
rect 590110 29574 590730 29658
rect 590110 29338 590142 29574
rect 590378 29338 590462 29574
rect 590698 29338 590730 29574
rect 590110 -5146 590730 29338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 693614 591690 710042
rect 591070 693378 591102 693614
rect 591338 693378 591422 693614
rect 591658 693378 591690 693614
rect 591070 693294 591690 693378
rect 591070 693058 591102 693294
rect 591338 693058 591422 693294
rect 591658 693058 591690 693294
rect 591070 653614 591690 693058
rect 591070 653378 591102 653614
rect 591338 653378 591422 653614
rect 591658 653378 591690 653614
rect 591070 653294 591690 653378
rect 591070 653058 591102 653294
rect 591338 653058 591422 653294
rect 591658 653058 591690 653294
rect 591070 613614 591690 653058
rect 591070 613378 591102 613614
rect 591338 613378 591422 613614
rect 591658 613378 591690 613614
rect 591070 613294 591690 613378
rect 591070 613058 591102 613294
rect 591338 613058 591422 613294
rect 591658 613058 591690 613294
rect 591070 573614 591690 613058
rect 591070 573378 591102 573614
rect 591338 573378 591422 573614
rect 591658 573378 591690 573614
rect 591070 573294 591690 573378
rect 591070 573058 591102 573294
rect 591338 573058 591422 573294
rect 591658 573058 591690 573294
rect 591070 533614 591690 573058
rect 591070 533378 591102 533614
rect 591338 533378 591422 533614
rect 591658 533378 591690 533614
rect 591070 533294 591690 533378
rect 591070 533058 591102 533294
rect 591338 533058 591422 533294
rect 591658 533058 591690 533294
rect 591070 493614 591690 533058
rect 591070 493378 591102 493614
rect 591338 493378 591422 493614
rect 591658 493378 591690 493614
rect 591070 493294 591690 493378
rect 591070 493058 591102 493294
rect 591338 493058 591422 493294
rect 591658 493058 591690 493294
rect 591070 453614 591690 493058
rect 591070 453378 591102 453614
rect 591338 453378 591422 453614
rect 591658 453378 591690 453614
rect 591070 453294 591690 453378
rect 591070 453058 591102 453294
rect 591338 453058 591422 453294
rect 591658 453058 591690 453294
rect 591070 413614 591690 453058
rect 591070 413378 591102 413614
rect 591338 413378 591422 413614
rect 591658 413378 591690 413614
rect 591070 413294 591690 413378
rect 591070 413058 591102 413294
rect 591338 413058 591422 413294
rect 591658 413058 591690 413294
rect 591070 373614 591690 413058
rect 591070 373378 591102 373614
rect 591338 373378 591422 373614
rect 591658 373378 591690 373614
rect 591070 373294 591690 373378
rect 591070 373058 591102 373294
rect 591338 373058 591422 373294
rect 591658 373058 591690 373294
rect 591070 333614 591690 373058
rect 591070 333378 591102 333614
rect 591338 333378 591422 333614
rect 591658 333378 591690 333614
rect 591070 333294 591690 333378
rect 591070 333058 591102 333294
rect 591338 333058 591422 333294
rect 591658 333058 591690 333294
rect 591070 293614 591690 333058
rect 591070 293378 591102 293614
rect 591338 293378 591422 293614
rect 591658 293378 591690 293614
rect 591070 293294 591690 293378
rect 591070 293058 591102 293294
rect 591338 293058 591422 293294
rect 591658 293058 591690 293294
rect 591070 253614 591690 293058
rect 591070 253378 591102 253614
rect 591338 253378 591422 253614
rect 591658 253378 591690 253614
rect 591070 253294 591690 253378
rect 591070 253058 591102 253294
rect 591338 253058 591422 253294
rect 591658 253058 591690 253294
rect 591070 213614 591690 253058
rect 591070 213378 591102 213614
rect 591338 213378 591422 213614
rect 591658 213378 591690 213614
rect 591070 213294 591690 213378
rect 591070 213058 591102 213294
rect 591338 213058 591422 213294
rect 591658 213058 591690 213294
rect 591070 173614 591690 213058
rect 591070 173378 591102 173614
rect 591338 173378 591422 173614
rect 591658 173378 591690 173614
rect 591070 173294 591690 173378
rect 591070 173058 591102 173294
rect 591338 173058 591422 173294
rect 591658 173058 591690 173294
rect 591070 133614 591690 173058
rect 591070 133378 591102 133614
rect 591338 133378 591422 133614
rect 591658 133378 591690 133614
rect 591070 133294 591690 133378
rect 591070 133058 591102 133294
rect 591338 133058 591422 133294
rect 591658 133058 591690 133294
rect 591070 93614 591690 133058
rect 591070 93378 591102 93614
rect 591338 93378 591422 93614
rect 591658 93378 591690 93614
rect 591070 93294 591690 93378
rect 591070 93058 591102 93294
rect 591338 93058 591422 93294
rect 591658 93058 591690 93294
rect 591070 53614 591690 93058
rect 591070 53378 591102 53614
rect 591338 53378 591422 53614
rect 591658 53378 591690 53614
rect 591070 53294 591690 53378
rect 591070 53058 591102 53294
rect 591338 53058 591422 53294
rect 591658 53058 591690 53294
rect 591070 13614 591690 53058
rect 591070 13378 591102 13614
rect 591338 13378 591422 13614
rect 591658 13378 591690 13614
rect 591070 13294 591690 13378
rect 591070 13058 591102 13294
rect 591338 13058 591422 13294
rect 591658 13058 591690 13294
rect 571954 -6342 571986 -6106
rect 572222 -6342 572306 -6106
rect 572542 -6342 572574 -6106
rect 571954 -6426 572574 -6342
rect 571954 -6662 571986 -6426
rect 572222 -6662 572306 -6426
rect 572542 -6662 572574 -6426
rect 571954 -7654 572574 -6662
rect 591070 -6106 591690 13058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 673614 592650 711002
rect 592030 673378 592062 673614
rect 592298 673378 592382 673614
rect 592618 673378 592650 673614
rect 592030 673294 592650 673378
rect 592030 673058 592062 673294
rect 592298 673058 592382 673294
rect 592618 673058 592650 673294
rect 592030 633614 592650 673058
rect 592030 633378 592062 633614
rect 592298 633378 592382 633614
rect 592618 633378 592650 633614
rect 592030 633294 592650 633378
rect 592030 633058 592062 633294
rect 592298 633058 592382 633294
rect 592618 633058 592650 633294
rect 592030 593614 592650 633058
rect 592030 593378 592062 593614
rect 592298 593378 592382 593614
rect 592618 593378 592650 593614
rect 592030 593294 592650 593378
rect 592030 593058 592062 593294
rect 592298 593058 592382 593294
rect 592618 593058 592650 593294
rect 592030 553614 592650 593058
rect 592030 553378 592062 553614
rect 592298 553378 592382 553614
rect 592618 553378 592650 553614
rect 592030 553294 592650 553378
rect 592030 553058 592062 553294
rect 592298 553058 592382 553294
rect 592618 553058 592650 553294
rect 592030 513614 592650 553058
rect 592030 513378 592062 513614
rect 592298 513378 592382 513614
rect 592618 513378 592650 513614
rect 592030 513294 592650 513378
rect 592030 513058 592062 513294
rect 592298 513058 592382 513294
rect 592618 513058 592650 513294
rect 592030 473614 592650 513058
rect 592030 473378 592062 473614
rect 592298 473378 592382 473614
rect 592618 473378 592650 473614
rect 592030 473294 592650 473378
rect 592030 473058 592062 473294
rect 592298 473058 592382 473294
rect 592618 473058 592650 473294
rect 592030 433614 592650 473058
rect 592030 433378 592062 433614
rect 592298 433378 592382 433614
rect 592618 433378 592650 433614
rect 592030 433294 592650 433378
rect 592030 433058 592062 433294
rect 592298 433058 592382 433294
rect 592618 433058 592650 433294
rect 592030 393614 592650 433058
rect 592030 393378 592062 393614
rect 592298 393378 592382 393614
rect 592618 393378 592650 393614
rect 592030 393294 592650 393378
rect 592030 393058 592062 393294
rect 592298 393058 592382 393294
rect 592618 393058 592650 393294
rect 592030 353614 592650 393058
rect 592030 353378 592062 353614
rect 592298 353378 592382 353614
rect 592618 353378 592650 353614
rect 592030 353294 592650 353378
rect 592030 353058 592062 353294
rect 592298 353058 592382 353294
rect 592618 353058 592650 353294
rect 592030 313614 592650 353058
rect 592030 313378 592062 313614
rect 592298 313378 592382 313614
rect 592618 313378 592650 313614
rect 592030 313294 592650 313378
rect 592030 313058 592062 313294
rect 592298 313058 592382 313294
rect 592618 313058 592650 313294
rect 592030 273614 592650 313058
rect 592030 273378 592062 273614
rect 592298 273378 592382 273614
rect 592618 273378 592650 273614
rect 592030 273294 592650 273378
rect 592030 273058 592062 273294
rect 592298 273058 592382 273294
rect 592618 273058 592650 273294
rect 592030 233614 592650 273058
rect 592030 233378 592062 233614
rect 592298 233378 592382 233614
rect 592618 233378 592650 233614
rect 592030 233294 592650 233378
rect 592030 233058 592062 233294
rect 592298 233058 592382 233294
rect 592618 233058 592650 233294
rect 592030 193614 592650 233058
rect 592030 193378 592062 193614
rect 592298 193378 592382 193614
rect 592618 193378 592650 193614
rect 592030 193294 592650 193378
rect 592030 193058 592062 193294
rect 592298 193058 592382 193294
rect 592618 193058 592650 193294
rect 592030 153614 592650 193058
rect 592030 153378 592062 153614
rect 592298 153378 592382 153614
rect 592618 153378 592650 153614
rect 592030 153294 592650 153378
rect 592030 153058 592062 153294
rect 592298 153058 592382 153294
rect 592618 153058 592650 153294
rect 592030 113614 592650 153058
rect 592030 113378 592062 113614
rect 592298 113378 592382 113614
rect 592618 113378 592650 113614
rect 592030 113294 592650 113378
rect 592030 113058 592062 113294
rect 592298 113058 592382 113294
rect 592618 113058 592650 113294
rect 592030 73614 592650 113058
rect 592030 73378 592062 73614
rect 592298 73378 592382 73614
rect 592618 73378 592650 73614
rect 592030 73294 592650 73378
rect 592030 73058 592062 73294
rect 592298 73058 592382 73294
rect 592618 73058 592650 73294
rect 592030 33614 592650 73058
rect 592030 33378 592062 33614
rect 592298 33378 592382 33614
rect 592618 33378 592650 33614
rect 592030 33294 592650 33378
rect 592030 33058 592062 33294
rect 592298 33058 592382 33294
rect 592618 33058 592650 33294
rect 592030 -7066 592650 33058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 673378 -8458 673614
rect -8374 673378 -8138 673614
rect -8694 673058 -8458 673294
rect -8374 673058 -8138 673294
rect -8694 633378 -8458 633614
rect -8374 633378 -8138 633614
rect -8694 633058 -8458 633294
rect -8374 633058 -8138 633294
rect -8694 593378 -8458 593614
rect -8374 593378 -8138 593614
rect -8694 593058 -8458 593294
rect -8374 593058 -8138 593294
rect -8694 553378 -8458 553614
rect -8374 553378 -8138 553614
rect -8694 553058 -8458 553294
rect -8374 553058 -8138 553294
rect -8694 513378 -8458 513614
rect -8374 513378 -8138 513614
rect -8694 513058 -8458 513294
rect -8374 513058 -8138 513294
rect -8694 473378 -8458 473614
rect -8374 473378 -8138 473614
rect -8694 473058 -8458 473294
rect -8374 473058 -8138 473294
rect -8694 433378 -8458 433614
rect -8374 433378 -8138 433614
rect -8694 433058 -8458 433294
rect -8374 433058 -8138 433294
rect -8694 393378 -8458 393614
rect -8374 393378 -8138 393614
rect -8694 393058 -8458 393294
rect -8374 393058 -8138 393294
rect -8694 353378 -8458 353614
rect -8374 353378 -8138 353614
rect -8694 353058 -8458 353294
rect -8374 353058 -8138 353294
rect -8694 313378 -8458 313614
rect -8374 313378 -8138 313614
rect -8694 313058 -8458 313294
rect -8374 313058 -8138 313294
rect -8694 273378 -8458 273614
rect -8374 273378 -8138 273614
rect -8694 273058 -8458 273294
rect -8374 273058 -8138 273294
rect -8694 233378 -8458 233614
rect -8374 233378 -8138 233614
rect -8694 233058 -8458 233294
rect -8374 233058 -8138 233294
rect -8694 193378 -8458 193614
rect -8374 193378 -8138 193614
rect -8694 193058 -8458 193294
rect -8374 193058 -8138 193294
rect -8694 153378 -8458 153614
rect -8374 153378 -8138 153614
rect -8694 153058 -8458 153294
rect -8374 153058 -8138 153294
rect -8694 113378 -8458 113614
rect -8374 113378 -8138 113614
rect -8694 113058 -8458 113294
rect -8374 113058 -8138 113294
rect -8694 73378 -8458 73614
rect -8374 73378 -8138 73614
rect -8694 73058 -8458 73294
rect -8374 73058 -8138 73294
rect -8694 33378 -8458 33614
rect -8374 33378 -8138 33614
rect -8694 33058 -8458 33294
rect -8374 33058 -8138 33294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 11986 710362 12222 710598
rect 12306 710362 12542 710598
rect 11986 710042 12222 710278
rect 12306 710042 12542 710278
rect -7734 693378 -7498 693614
rect -7414 693378 -7178 693614
rect -7734 693058 -7498 693294
rect -7414 693058 -7178 693294
rect -7734 653378 -7498 653614
rect -7414 653378 -7178 653614
rect -7734 653058 -7498 653294
rect -7414 653058 -7178 653294
rect -7734 613378 -7498 613614
rect -7414 613378 -7178 613614
rect -7734 613058 -7498 613294
rect -7414 613058 -7178 613294
rect -7734 573378 -7498 573614
rect -7414 573378 -7178 573614
rect -7734 573058 -7498 573294
rect -7414 573058 -7178 573294
rect -7734 533378 -7498 533614
rect -7414 533378 -7178 533614
rect -7734 533058 -7498 533294
rect -7414 533058 -7178 533294
rect -7734 493378 -7498 493614
rect -7414 493378 -7178 493614
rect -7734 493058 -7498 493294
rect -7414 493058 -7178 493294
rect -7734 453378 -7498 453614
rect -7414 453378 -7178 453614
rect -7734 453058 -7498 453294
rect -7414 453058 -7178 453294
rect -7734 413378 -7498 413614
rect -7414 413378 -7178 413614
rect -7734 413058 -7498 413294
rect -7414 413058 -7178 413294
rect -7734 373378 -7498 373614
rect -7414 373378 -7178 373614
rect -7734 373058 -7498 373294
rect -7414 373058 -7178 373294
rect -7734 333378 -7498 333614
rect -7414 333378 -7178 333614
rect -7734 333058 -7498 333294
rect -7414 333058 -7178 333294
rect -7734 293378 -7498 293614
rect -7414 293378 -7178 293614
rect -7734 293058 -7498 293294
rect -7414 293058 -7178 293294
rect -7734 253378 -7498 253614
rect -7414 253378 -7178 253614
rect -7734 253058 -7498 253294
rect -7414 253058 -7178 253294
rect -7734 213378 -7498 213614
rect -7414 213378 -7178 213614
rect -7734 213058 -7498 213294
rect -7414 213058 -7178 213294
rect -7734 173378 -7498 173614
rect -7414 173378 -7178 173614
rect -7734 173058 -7498 173294
rect -7414 173058 -7178 173294
rect -7734 133378 -7498 133614
rect -7414 133378 -7178 133614
rect -7734 133058 -7498 133294
rect -7414 133058 -7178 133294
rect -7734 93378 -7498 93614
rect -7414 93378 -7178 93614
rect -7734 93058 -7498 93294
rect -7414 93058 -7178 93294
rect -7734 53378 -7498 53614
rect -7414 53378 -7178 53614
rect -7734 53058 -7498 53294
rect -7414 53058 -7178 53294
rect -7734 13378 -7498 13614
rect -7414 13378 -7178 13614
rect -7734 13058 -7498 13294
rect -7414 13058 -7178 13294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669658 -6538 669894
rect -6454 669658 -6218 669894
rect -6774 669338 -6538 669574
rect -6454 669338 -6218 669574
rect -6774 629658 -6538 629894
rect -6454 629658 -6218 629894
rect -6774 629338 -6538 629574
rect -6454 629338 -6218 629574
rect -6774 589658 -6538 589894
rect -6454 589658 -6218 589894
rect -6774 589338 -6538 589574
rect -6454 589338 -6218 589574
rect -6774 549658 -6538 549894
rect -6454 549658 -6218 549894
rect -6774 549338 -6538 549574
rect -6454 549338 -6218 549574
rect -6774 509658 -6538 509894
rect -6454 509658 -6218 509894
rect -6774 509338 -6538 509574
rect -6454 509338 -6218 509574
rect -6774 469658 -6538 469894
rect -6454 469658 -6218 469894
rect -6774 469338 -6538 469574
rect -6454 469338 -6218 469574
rect -6774 429658 -6538 429894
rect -6454 429658 -6218 429894
rect -6774 429338 -6538 429574
rect -6454 429338 -6218 429574
rect -6774 389658 -6538 389894
rect -6454 389658 -6218 389894
rect -6774 389338 -6538 389574
rect -6454 389338 -6218 389574
rect -6774 349658 -6538 349894
rect -6454 349658 -6218 349894
rect -6774 349338 -6538 349574
rect -6454 349338 -6218 349574
rect -6774 309658 -6538 309894
rect -6454 309658 -6218 309894
rect -6774 309338 -6538 309574
rect -6454 309338 -6218 309574
rect -6774 269658 -6538 269894
rect -6454 269658 -6218 269894
rect -6774 269338 -6538 269574
rect -6454 269338 -6218 269574
rect -6774 229658 -6538 229894
rect -6454 229658 -6218 229894
rect -6774 229338 -6538 229574
rect -6454 229338 -6218 229574
rect -6774 189658 -6538 189894
rect -6454 189658 -6218 189894
rect -6774 189338 -6538 189574
rect -6454 189338 -6218 189574
rect -6774 149658 -6538 149894
rect -6454 149658 -6218 149894
rect -6774 149338 -6538 149574
rect -6454 149338 -6218 149574
rect -6774 109658 -6538 109894
rect -6454 109658 -6218 109894
rect -6774 109338 -6538 109574
rect -6454 109338 -6218 109574
rect -6774 69658 -6538 69894
rect -6454 69658 -6218 69894
rect -6774 69338 -6538 69574
rect -6454 69338 -6218 69574
rect -6774 29658 -6538 29894
rect -6454 29658 -6218 29894
rect -6774 29338 -6538 29574
rect -6454 29338 -6218 29574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 8266 708442 8502 708678
rect 8586 708442 8822 708678
rect 8266 708122 8502 708358
rect 8586 708122 8822 708358
rect -5814 689658 -5578 689894
rect -5494 689658 -5258 689894
rect -5814 689338 -5578 689574
rect -5494 689338 -5258 689574
rect -5814 649658 -5578 649894
rect -5494 649658 -5258 649894
rect -5814 649338 -5578 649574
rect -5494 649338 -5258 649574
rect -5814 609658 -5578 609894
rect -5494 609658 -5258 609894
rect -5814 609338 -5578 609574
rect -5494 609338 -5258 609574
rect -5814 569658 -5578 569894
rect -5494 569658 -5258 569894
rect -5814 569338 -5578 569574
rect -5494 569338 -5258 569574
rect -5814 529658 -5578 529894
rect -5494 529658 -5258 529894
rect -5814 529338 -5578 529574
rect -5494 529338 -5258 529574
rect -5814 489658 -5578 489894
rect -5494 489658 -5258 489894
rect -5814 489338 -5578 489574
rect -5494 489338 -5258 489574
rect -5814 449658 -5578 449894
rect -5494 449658 -5258 449894
rect -5814 449338 -5578 449574
rect -5494 449338 -5258 449574
rect -5814 409658 -5578 409894
rect -5494 409658 -5258 409894
rect -5814 409338 -5578 409574
rect -5494 409338 -5258 409574
rect -5814 369658 -5578 369894
rect -5494 369658 -5258 369894
rect -5814 369338 -5578 369574
rect -5494 369338 -5258 369574
rect -5814 329658 -5578 329894
rect -5494 329658 -5258 329894
rect -5814 329338 -5578 329574
rect -5494 329338 -5258 329574
rect -5814 289658 -5578 289894
rect -5494 289658 -5258 289894
rect -5814 289338 -5578 289574
rect -5494 289338 -5258 289574
rect -5814 249658 -5578 249894
rect -5494 249658 -5258 249894
rect -5814 249338 -5578 249574
rect -5494 249338 -5258 249574
rect -5814 209658 -5578 209894
rect -5494 209658 -5258 209894
rect -5814 209338 -5578 209574
rect -5494 209338 -5258 209574
rect -5814 169658 -5578 169894
rect -5494 169658 -5258 169894
rect -5814 169338 -5578 169574
rect -5494 169338 -5258 169574
rect -5814 129658 -5578 129894
rect -5494 129658 -5258 129894
rect -5814 129338 -5578 129574
rect -5494 129338 -5258 129574
rect -5814 89658 -5578 89894
rect -5494 89658 -5258 89894
rect -5814 89338 -5578 89574
rect -5494 89338 -5258 89574
rect -5814 49658 -5578 49894
rect -5494 49658 -5258 49894
rect -5814 49338 -5578 49574
rect -5494 49338 -5258 49574
rect -5814 9658 -5578 9894
rect -5494 9658 -5258 9894
rect -5814 9338 -5578 9574
rect -5494 9338 -5258 9574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 665938 -4618 666174
rect -4534 665938 -4298 666174
rect -4854 665618 -4618 665854
rect -4534 665618 -4298 665854
rect -4854 625938 -4618 626174
rect -4534 625938 -4298 626174
rect -4854 625618 -4618 625854
rect -4534 625618 -4298 625854
rect -4854 585938 -4618 586174
rect -4534 585938 -4298 586174
rect -4854 585618 -4618 585854
rect -4534 585618 -4298 585854
rect -4854 545938 -4618 546174
rect -4534 545938 -4298 546174
rect -4854 545618 -4618 545854
rect -4534 545618 -4298 545854
rect -4854 505938 -4618 506174
rect -4534 505938 -4298 506174
rect -4854 505618 -4618 505854
rect -4534 505618 -4298 505854
rect -4854 465938 -4618 466174
rect -4534 465938 -4298 466174
rect -4854 465618 -4618 465854
rect -4534 465618 -4298 465854
rect -4854 425938 -4618 426174
rect -4534 425938 -4298 426174
rect -4854 425618 -4618 425854
rect -4534 425618 -4298 425854
rect -4854 385938 -4618 386174
rect -4534 385938 -4298 386174
rect -4854 385618 -4618 385854
rect -4534 385618 -4298 385854
rect -4854 345938 -4618 346174
rect -4534 345938 -4298 346174
rect -4854 345618 -4618 345854
rect -4534 345618 -4298 345854
rect -4854 305938 -4618 306174
rect -4534 305938 -4298 306174
rect -4854 305618 -4618 305854
rect -4534 305618 -4298 305854
rect -4854 265938 -4618 266174
rect -4534 265938 -4298 266174
rect -4854 265618 -4618 265854
rect -4534 265618 -4298 265854
rect -4854 225938 -4618 226174
rect -4534 225938 -4298 226174
rect -4854 225618 -4618 225854
rect -4534 225618 -4298 225854
rect -4854 185938 -4618 186174
rect -4534 185938 -4298 186174
rect -4854 185618 -4618 185854
rect -4534 185618 -4298 185854
rect -4854 145938 -4618 146174
rect -4534 145938 -4298 146174
rect -4854 145618 -4618 145854
rect -4534 145618 -4298 145854
rect -4854 105938 -4618 106174
rect -4534 105938 -4298 106174
rect -4854 105618 -4618 105854
rect -4534 105618 -4298 105854
rect -4854 65938 -4618 66174
rect -4534 65938 -4298 66174
rect -4854 65618 -4618 65854
rect -4534 65618 -4298 65854
rect -4854 25938 -4618 26174
rect -4534 25938 -4298 26174
rect -4854 25618 -4618 25854
rect -4534 25618 -4298 25854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 4546 706522 4782 706758
rect 4866 706522 5102 706758
rect 4546 706202 4782 706438
rect 4866 706202 5102 706438
rect -3894 685938 -3658 686174
rect -3574 685938 -3338 686174
rect -3894 685618 -3658 685854
rect -3574 685618 -3338 685854
rect -3894 645938 -3658 646174
rect -3574 645938 -3338 646174
rect -3894 645618 -3658 645854
rect -3574 645618 -3338 645854
rect -3894 605938 -3658 606174
rect -3574 605938 -3338 606174
rect -3894 605618 -3658 605854
rect -3574 605618 -3338 605854
rect -3894 565938 -3658 566174
rect -3574 565938 -3338 566174
rect -3894 565618 -3658 565854
rect -3574 565618 -3338 565854
rect -3894 525938 -3658 526174
rect -3574 525938 -3338 526174
rect -3894 525618 -3658 525854
rect -3574 525618 -3338 525854
rect -3894 485938 -3658 486174
rect -3574 485938 -3338 486174
rect -3894 485618 -3658 485854
rect -3574 485618 -3338 485854
rect -3894 445938 -3658 446174
rect -3574 445938 -3338 446174
rect -3894 445618 -3658 445854
rect -3574 445618 -3338 445854
rect -3894 405938 -3658 406174
rect -3574 405938 -3338 406174
rect -3894 405618 -3658 405854
rect -3574 405618 -3338 405854
rect -3894 365938 -3658 366174
rect -3574 365938 -3338 366174
rect -3894 365618 -3658 365854
rect -3574 365618 -3338 365854
rect -3894 325938 -3658 326174
rect -3574 325938 -3338 326174
rect -3894 325618 -3658 325854
rect -3574 325618 -3338 325854
rect -3894 285938 -3658 286174
rect -3574 285938 -3338 286174
rect -3894 285618 -3658 285854
rect -3574 285618 -3338 285854
rect -3894 245938 -3658 246174
rect -3574 245938 -3338 246174
rect -3894 245618 -3658 245854
rect -3574 245618 -3338 245854
rect -3894 205938 -3658 206174
rect -3574 205938 -3338 206174
rect -3894 205618 -3658 205854
rect -3574 205618 -3338 205854
rect -3894 165938 -3658 166174
rect -3574 165938 -3338 166174
rect -3894 165618 -3658 165854
rect -3574 165618 -3338 165854
rect -3894 125938 -3658 126174
rect -3574 125938 -3338 126174
rect -3894 125618 -3658 125854
rect -3574 125618 -3338 125854
rect -3894 85938 -3658 86174
rect -3574 85938 -3338 86174
rect -3894 85618 -3658 85854
rect -3574 85618 -3338 85854
rect -3894 45938 -3658 46174
rect -3574 45938 -3338 46174
rect -3894 45618 -3658 45854
rect -3574 45618 -3338 45854
rect -3894 5938 -3658 6174
rect -3574 5938 -3338 6174
rect -3894 5618 -3658 5854
rect -3574 5618 -3338 5854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 662218 -2698 662454
rect -2614 662218 -2378 662454
rect -2934 661898 -2698 662134
rect -2614 661898 -2378 662134
rect -2934 622218 -2698 622454
rect -2614 622218 -2378 622454
rect -2934 621898 -2698 622134
rect -2614 621898 -2378 622134
rect -2934 582218 -2698 582454
rect -2614 582218 -2378 582454
rect -2934 581898 -2698 582134
rect -2614 581898 -2378 582134
rect -2934 542218 -2698 542454
rect -2614 542218 -2378 542454
rect -2934 541898 -2698 542134
rect -2614 541898 -2378 542134
rect -2934 502218 -2698 502454
rect -2614 502218 -2378 502454
rect -2934 501898 -2698 502134
rect -2614 501898 -2378 502134
rect -2934 462218 -2698 462454
rect -2614 462218 -2378 462454
rect -2934 461898 -2698 462134
rect -2614 461898 -2378 462134
rect -2934 422218 -2698 422454
rect -2614 422218 -2378 422454
rect -2934 421898 -2698 422134
rect -2614 421898 -2378 422134
rect -2934 382218 -2698 382454
rect -2614 382218 -2378 382454
rect -2934 381898 -2698 382134
rect -2614 381898 -2378 382134
rect -2934 342218 -2698 342454
rect -2614 342218 -2378 342454
rect -2934 341898 -2698 342134
rect -2614 341898 -2378 342134
rect -2934 302218 -2698 302454
rect -2614 302218 -2378 302454
rect -2934 301898 -2698 302134
rect -2614 301898 -2378 302134
rect -2934 262218 -2698 262454
rect -2614 262218 -2378 262454
rect -2934 261898 -2698 262134
rect -2614 261898 -2378 262134
rect -2934 222218 -2698 222454
rect -2614 222218 -2378 222454
rect -2934 221898 -2698 222134
rect -2614 221898 -2378 222134
rect -2934 182218 -2698 182454
rect -2614 182218 -2378 182454
rect -2934 181898 -2698 182134
rect -2614 181898 -2378 182134
rect -2934 142218 -2698 142454
rect -2614 142218 -2378 142454
rect -2934 141898 -2698 142134
rect -2614 141898 -2378 142134
rect -2934 102218 -2698 102454
rect -2614 102218 -2378 102454
rect -2934 101898 -2698 102134
rect -2614 101898 -2378 102134
rect -2934 62218 -2698 62454
rect -2614 62218 -2378 62454
rect -2934 61898 -2698 62134
rect -2614 61898 -2378 62134
rect -2934 22218 -2698 22454
rect -2614 22218 -2378 22454
rect -2934 21898 -2698 22134
rect -2614 21898 -2378 22134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 682218 -1738 682454
rect -1654 682218 -1418 682454
rect -1974 681898 -1738 682134
rect -1654 681898 -1418 682134
rect -1974 642218 -1738 642454
rect -1654 642218 -1418 642454
rect -1974 641898 -1738 642134
rect -1654 641898 -1418 642134
rect -1974 602218 -1738 602454
rect -1654 602218 -1418 602454
rect -1974 601898 -1738 602134
rect -1654 601898 -1418 602134
rect -1974 562218 -1738 562454
rect -1654 562218 -1418 562454
rect -1974 561898 -1738 562134
rect -1654 561898 -1418 562134
rect -1974 522218 -1738 522454
rect -1654 522218 -1418 522454
rect -1974 521898 -1738 522134
rect -1654 521898 -1418 522134
rect -1974 482218 -1738 482454
rect -1654 482218 -1418 482454
rect -1974 481898 -1738 482134
rect -1654 481898 -1418 482134
rect -1974 442218 -1738 442454
rect -1654 442218 -1418 442454
rect -1974 441898 -1738 442134
rect -1654 441898 -1418 442134
rect -1974 402218 -1738 402454
rect -1654 402218 -1418 402454
rect -1974 401898 -1738 402134
rect -1654 401898 -1418 402134
rect -1974 362218 -1738 362454
rect -1654 362218 -1418 362454
rect -1974 361898 -1738 362134
rect -1654 361898 -1418 362134
rect -1974 322218 -1738 322454
rect -1654 322218 -1418 322454
rect -1974 321898 -1738 322134
rect -1654 321898 -1418 322134
rect -1974 282218 -1738 282454
rect -1654 282218 -1418 282454
rect -1974 281898 -1738 282134
rect -1654 281898 -1418 282134
rect -1974 242218 -1738 242454
rect -1654 242218 -1418 242454
rect -1974 241898 -1738 242134
rect -1654 241898 -1418 242134
rect -1974 202218 -1738 202454
rect -1654 202218 -1418 202454
rect -1974 201898 -1738 202134
rect -1654 201898 -1418 202134
rect -1974 162218 -1738 162454
rect -1654 162218 -1418 162454
rect -1974 161898 -1738 162134
rect -1654 161898 -1418 162134
rect -1974 122218 -1738 122454
rect -1654 122218 -1418 122454
rect -1974 121898 -1738 122134
rect -1654 121898 -1418 122134
rect -1974 82218 -1738 82454
rect -1654 82218 -1418 82454
rect -1974 81898 -1738 82134
rect -1654 81898 -1418 82134
rect -1974 42218 -1738 42454
rect -1654 42218 -1418 42454
rect -1974 41898 -1738 42134
rect -1654 41898 -1418 42134
rect -1974 2218 -1738 2454
rect -1654 2218 -1418 2454
rect -1974 1898 -1738 2134
rect -1654 1898 -1418 2134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 826 704602 1062 704838
rect 1146 704602 1382 704838
rect 826 704282 1062 704518
rect 1146 704282 1382 704518
rect 826 682218 1062 682454
rect 1146 682218 1382 682454
rect 826 681898 1062 682134
rect 1146 681898 1382 682134
rect 826 642218 1062 642454
rect 1146 642218 1382 642454
rect 826 641898 1062 642134
rect 1146 641898 1382 642134
rect 826 602218 1062 602454
rect 1146 602218 1382 602454
rect 826 601898 1062 602134
rect 1146 601898 1382 602134
rect 826 562218 1062 562454
rect 1146 562218 1382 562454
rect 826 561898 1062 562134
rect 1146 561898 1382 562134
rect 826 522218 1062 522454
rect 1146 522218 1382 522454
rect 826 521898 1062 522134
rect 1146 521898 1382 522134
rect 826 482218 1062 482454
rect 1146 482218 1382 482454
rect 826 481898 1062 482134
rect 1146 481898 1382 482134
rect 826 442218 1062 442454
rect 1146 442218 1382 442454
rect 826 441898 1062 442134
rect 1146 441898 1382 442134
rect 826 402218 1062 402454
rect 1146 402218 1382 402454
rect 826 401898 1062 402134
rect 1146 401898 1382 402134
rect 826 362218 1062 362454
rect 1146 362218 1382 362454
rect 826 361898 1062 362134
rect 1146 361898 1382 362134
rect 826 322218 1062 322454
rect 1146 322218 1382 322454
rect 826 321898 1062 322134
rect 1146 321898 1382 322134
rect 826 282218 1062 282454
rect 1146 282218 1382 282454
rect 826 281898 1062 282134
rect 1146 281898 1382 282134
rect 826 242218 1062 242454
rect 1146 242218 1382 242454
rect 826 241898 1062 242134
rect 1146 241898 1382 242134
rect 826 202218 1062 202454
rect 1146 202218 1382 202454
rect 826 201898 1062 202134
rect 1146 201898 1382 202134
rect 826 162218 1062 162454
rect 1146 162218 1382 162454
rect 826 161898 1062 162134
rect 1146 161898 1382 162134
rect 826 122218 1062 122454
rect 1146 122218 1382 122454
rect 826 121898 1062 122134
rect 1146 121898 1382 122134
rect 826 82218 1062 82454
rect 1146 82218 1382 82454
rect 826 81898 1062 82134
rect 1146 81898 1382 82134
rect 826 42218 1062 42454
rect 1146 42218 1382 42454
rect 826 41898 1062 42134
rect 1146 41898 1382 42134
rect 826 2218 1062 2454
rect 1146 2218 1382 2454
rect 826 1898 1062 2134
rect 1146 1898 1382 2134
rect 826 -582 1062 -346
rect 1146 -582 1382 -346
rect 826 -902 1062 -666
rect 1146 -902 1382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 4546 685938 4782 686174
rect 4866 685938 5102 686174
rect 4546 685618 4782 685854
rect 4866 685618 5102 685854
rect 4546 645938 4782 646174
rect 4866 645938 5102 646174
rect 4546 645618 4782 645854
rect 4866 645618 5102 645854
rect 4546 605938 4782 606174
rect 4866 605938 5102 606174
rect 4546 605618 4782 605854
rect 4866 605618 5102 605854
rect 4546 565938 4782 566174
rect 4866 565938 5102 566174
rect 4546 565618 4782 565854
rect 4866 565618 5102 565854
rect 4546 525938 4782 526174
rect 4866 525938 5102 526174
rect 4546 525618 4782 525854
rect 4866 525618 5102 525854
rect 4546 485938 4782 486174
rect 4866 485938 5102 486174
rect 4546 485618 4782 485854
rect 4866 485618 5102 485854
rect 4546 445938 4782 446174
rect 4866 445938 5102 446174
rect 4546 445618 4782 445854
rect 4866 445618 5102 445854
rect 4546 405938 4782 406174
rect 4866 405938 5102 406174
rect 4546 405618 4782 405854
rect 4866 405618 5102 405854
rect 4546 365938 4782 366174
rect 4866 365938 5102 366174
rect 4546 365618 4782 365854
rect 4866 365618 5102 365854
rect 4546 325938 4782 326174
rect 4866 325938 5102 326174
rect 4546 325618 4782 325854
rect 4866 325618 5102 325854
rect 4546 285938 4782 286174
rect 4866 285938 5102 286174
rect 4546 285618 4782 285854
rect 4866 285618 5102 285854
rect 4546 245938 4782 246174
rect 4866 245938 5102 246174
rect 4546 245618 4782 245854
rect 4866 245618 5102 245854
rect 4546 205938 4782 206174
rect 4866 205938 5102 206174
rect 4546 205618 4782 205854
rect 4866 205618 5102 205854
rect 4546 165938 4782 166174
rect 4866 165938 5102 166174
rect 4546 165618 4782 165854
rect 4866 165618 5102 165854
rect 4546 125938 4782 126174
rect 4866 125938 5102 126174
rect 4546 125618 4782 125854
rect 4866 125618 5102 125854
rect 4546 85938 4782 86174
rect 4866 85938 5102 86174
rect 4546 85618 4782 85854
rect 4866 85618 5102 85854
rect 4546 45938 4782 46174
rect 4866 45938 5102 46174
rect 4546 45618 4782 45854
rect 4866 45618 5102 45854
rect 4546 5938 4782 6174
rect 4866 5938 5102 6174
rect 4546 5618 4782 5854
rect 4866 5618 5102 5854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 4546 -2502 4782 -2266
rect 4866 -2502 5102 -2266
rect 4546 -2822 4782 -2586
rect 4866 -2822 5102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 8266 689658 8502 689894
rect 8586 689658 8822 689894
rect 8266 689338 8502 689574
rect 8586 689338 8822 689574
rect 8266 649658 8502 649894
rect 8586 649658 8822 649894
rect 8266 649338 8502 649574
rect 8586 649338 8822 649574
rect 8266 609658 8502 609894
rect 8586 609658 8822 609894
rect 8266 609338 8502 609574
rect 8586 609338 8822 609574
rect 8266 569658 8502 569894
rect 8586 569658 8822 569894
rect 8266 569338 8502 569574
rect 8586 569338 8822 569574
rect 8266 529658 8502 529894
rect 8586 529658 8822 529894
rect 8266 529338 8502 529574
rect 8586 529338 8822 529574
rect 8266 489658 8502 489894
rect 8586 489658 8822 489894
rect 8266 489338 8502 489574
rect 8586 489338 8822 489574
rect 8266 449658 8502 449894
rect 8586 449658 8822 449894
rect 8266 449338 8502 449574
rect 8586 449338 8822 449574
rect 8266 409658 8502 409894
rect 8586 409658 8822 409894
rect 8266 409338 8502 409574
rect 8586 409338 8822 409574
rect 8266 369658 8502 369894
rect 8586 369658 8822 369894
rect 8266 369338 8502 369574
rect 8586 369338 8822 369574
rect 8266 329658 8502 329894
rect 8586 329658 8822 329894
rect 8266 329338 8502 329574
rect 8586 329338 8822 329574
rect 8266 289658 8502 289894
rect 8586 289658 8822 289894
rect 8266 289338 8502 289574
rect 8586 289338 8822 289574
rect 8266 249658 8502 249894
rect 8586 249658 8822 249894
rect 8266 249338 8502 249574
rect 8586 249338 8822 249574
rect 8266 209658 8502 209894
rect 8586 209658 8822 209894
rect 8266 209338 8502 209574
rect 8586 209338 8822 209574
rect 8266 169658 8502 169894
rect 8586 169658 8822 169894
rect 8266 169338 8502 169574
rect 8586 169338 8822 169574
rect 8266 129658 8502 129894
rect 8586 129658 8822 129894
rect 8266 129338 8502 129574
rect 8586 129338 8822 129574
rect 8266 89658 8502 89894
rect 8586 89658 8822 89894
rect 8266 89338 8502 89574
rect 8586 89338 8822 89574
rect 8266 49658 8502 49894
rect 8586 49658 8822 49894
rect 8266 49338 8502 49574
rect 8586 49338 8822 49574
rect 8266 9658 8502 9894
rect 8586 9658 8822 9894
rect 8266 9338 8502 9574
rect 8586 9338 8822 9574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 8266 -4422 8502 -4186
rect 8586 -4422 8822 -4186
rect 8266 -4742 8502 -4506
rect 8586 -4742 8822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 31986 711322 32222 711558
rect 32306 711322 32542 711558
rect 31986 711002 32222 711238
rect 32306 711002 32542 711238
rect 28266 709402 28502 709638
rect 28586 709402 28822 709638
rect 28266 709082 28502 709318
rect 28586 709082 28822 709318
rect 24546 707482 24782 707718
rect 24866 707482 25102 707718
rect 24546 707162 24782 707398
rect 24866 707162 25102 707398
rect 11986 693378 12222 693614
rect 12306 693378 12542 693614
rect 11986 693058 12222 693294
rect 12306 693058 12542 693294
rect 11986 653378 12222 653614
rect 12306 653378 12542 653614
rect 11986 653058 12222 653294
rect 12306 653058 12542 653294
rect 11986 613378 12222 613614
rect 12306 613378 12542 613614
rect 11986 613058 12222 613294
rect 12306 613058 12542 613294
rect 11986 573378 12222 573614
rect 12306 573378 12542 573614
rect 11986 573058 12222 573294
rect 12306 573058 12542 573294
rect 11986 533378 12222 533614
rect 12306 533378 12542 533614
rect 11986 533058 12222 533294
rect 12306 533058 12542 533294
rect 11986 493378 12222 493614
rect 12306 493378 12542 493614
rect 11986 493058 12222 493294
rect 12306 493058 12542 493294
rect 11986 453378 12222 453614
rect 12306 453378 12542 453614
rect 11986 453058 12222 453294
rect 12306 453058 12542 453294
rect 11986 413378 12222 413614
rect 12306 413378 12542 413614
rect 11986 413058 12222 413294
rect 12306 413058 12542 413294
rect 11986 373378 12222 373614
rect 12306 373378 12542 373614
rect 11986 373058 12222 373294
rect 12306 373058 12542 373294
rect 11986 333378 12222 333614
rect 12306 333378 12542 333614
rect 11986 333058 12222 333294
rect 12306 333058 12542 333294
rect 11986 293378 12222 293614
rect 12306 293378 12542 293614
rect 11986 293058 12222 293294
rect 12306 293058 12542 293294
rect 11986 253378 12222 253614
rect 12306 253378 12542 253614
rect 11986 253058 12222 253294
rect 12306 253058 12542 253294
rect 11986 213378 12222 213614
rect 12306 213378 12542 213614
rect 11986 213058 12222 213294
rect 12306 213058 12542 213294
rect 11986 173378 12222 173614
rect 12306 173378 12542 173614
rect 11986 173058 12222 173294
rect 12306 173058 12542 173294
rect 11986 133378 12222 133614
rect 12306 133378 12542 133614
rect 11986 133058 12222 133294
rect 12306 133058 12542 133294
rect 11986 93378 12222 93614
rect 12306 93378 12542 93614
rect 11986 93058 12222 93294
rect 12306 93058 12542 93294
rect 11986 53378 12222 53614
rect 12306 53378 12542 53614
rect 11986 53058 12222 53294
rect 12306 53058 12542 53294
rect 11986 13378 12222 13614
rect 12306 13378 12542 13614
rect 11986 13058 12222 13294
rect 12306 13058 12542 13294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 20826 705562 21062 705798
rect 21146 705562 21382 705798
rect 20826 705242 21062 705478
rect 21146 705242 21382 705478
rect 20826 662218 21062 662454
rect 21146 662218 21382 662454
rect 20826 661898 21062 662134
rect 21146 661898 21382 662134
rect 20826 622218 21062 622454
rect 21146 622218 21382 622454
rect 20826 621898 21062 622134
rect 21146 621898 21382 622134
rect 20826 582218 21062 582454
rect 21146 582218 21382 582454
rect 20826 581898 21062 582134
rect 21146 581898 21382 582134
rect 20826 542218 21062 542454
rect 21146 542218 21382 542454
rect 20826 541898 21062 542134
rect 21146 541898 21382 542134
rect 20826 502218 21062 502454
rect 21146 502218 21382 502454
rect 20826 501898 21062 502134
rect 21146 501898 21382 502134
rect 20826 462218 21062 462454
rect 21146 462218 21382 462454
rect 20826 461898 21062 462134
rect 21146 461898 21382 462134
rect 20826 422218 21062 422454
rect 21146 422218 21382 422454
rect 20826 421898 21062 422134
rect 21146 421898 21382 422134
rect 20826 382218 21062 382454
rect 21146 382218 21382 382454
rect 20826 381898 21062 382134
rect 21146 381898 21382 382134
rect 20826 342218 21062 342454
rect 21146 342218 21382 342454
rect 20826 341898 21062 342134
rect 21146 341898 21382 342134
rect 20826 302218 21062 302454
rect 21146 302218 21382 302454
rect 20826 301898 21062 302134
rect 21146 301898 21382 302134
rect 20826 262218 21062 262454
rect 21146 262218 21382 262454
rect 20826 261898 21062 262134
rect 21146 261898 21382 262134
rect 20826 222218 21062 222454
rect 21146 222218 21382 222454
rect 20826 221898 21062 222134
rect 21146 221898 21382 222134
rect 20826 182218 21062 182454
rect 21146 182218 21382 182454
rect 20826 181898 21062 182134
rect 21146 181898 21382 182134
rect 20826 142218 21062 142454
rect 21146 142218 21382 142454
rect 20826 141898 21062 142134
rect 21146 141898 21382 142134
rect 20826 102218 21062 102454
rect 21146 102218 21382 102454
rect 20826 101898 21062 102134
rect 21146 101898 21382 102134
rect 20826 62218 21062 62454
rect 21146 62218 21382 62454
rect 20826 61898 21062 62134
rect 21146 61898 21382 62134
rect 20826 22218 21062 22454
rect 21146 22218 21382 22454
rect 20826 21898 21062 22134
rect 21146 21898 21382 22134
rect 20826 -1542 21062 -1306
rect 21146 -1542 21382 -1306
rect 20826 -1862 21062 -1626
rect 21146 -1862 21382 -1626
rect 24546 665938 24782 666174
rect 24866 665938 25102 666174
rect 24546 665618 24782 665854
rect 24866 665618 25102 665854
rect 24546 625938 24782 626174
rect 24866 625938 25102 626174
rect 24546 625618 24782 625854
rect 24866 625618 25102 625854
rect 24546 585938 24782 586174
rect 24866 585938 25102 586174
rect 24546 585618 24782 585854
rect 24866 585618 25102 585854
rect 24546 545938 24782 546174
rect 24866 545938 25102 546174
rect 24546 545618 24782 545854
rect 24866 545618 25102 545854
rect 24546 505938 24782 506174
rect 24866 505938 25102 506174
rect 24546 505618 24782 505854
rect 24866 505618 25102 505854
rect 24546 465938 24782 466174
rect 24866 465938 25102 466174
rect 24546 465618 24782 465854
rect 24866 465618 25102 465854
rect 24546 425938 24782 426174
rect 24866 425938 25102 426174
rect 24546 425618 24782 425854
rect 24866 425618 25102 425854
rect 24546 385938 24782 386174
rect 24866 385938 25102 386174
rect 24546 385618 24782 385854
rect 24866 385618 25102 385854
rect 24546 345938 24782 346174
rect 24866 345938 25102 346174
rect 24546 345618 24782 345854
rect 24866 345618 25102 345854
rect 24546 305938 24782 306174
rect 24866 305938 25102 306174
rect 24546 305618 24782 305854
rect 24866 305618 25102 305854
rect 24546 265938 24782 266174
rect 24866 265938 25102 266174
rect 24546 265618 24782 265854
rect 24866 265618 25102 265854
rect 24546 225938 24782 226174
rect 24866 225938 25102 226174
rect 24546 225618 24782 225854
rect 24866 225618 25102 225854
rect 24546 185938 24782 186174
rect 24866 185938 25102 186174
rect 24546 185618 24782 185854
rect 24866 185618 25102 185854
rect 24546 145938 24782 146174
rect 24866 145938 25102 146174
rect 24546 145618 24782 145854
rect 24866 145618 25102 145854
rect 24546 105938 24782 106174
rect 24866 105938 25102 106174
rect 24546 105618 24782 105854
rect 24866 105618 25102 105854
rect 24546 65938 24782 66174
rect 24866 65938 25102 66174
rect 24546 65618 24782 65854
rect 24866 65618 25102 65854
rect 24546 25938 24782 26174
rect 24866 25938 25102 26174
rect 24546 25618 24782 25854
rect 24866 25618 25102 25854
rect 24546 -3462 24782 -3226
rect 24866 -3462 25102 -3226
rect 24546 -3782 24782 -3546
rect 24866 -3782 25102 -3546
rect 28266 669658 28502 669894
rect 28586 669658 28822 669894
rect 28266 669338 28502 669574
rect 28586 669338 28822 669574
rect 28266 629658 28502 629894
rect 28586 629658 28822 629894
rect 28266 629338 28502 629574
rect 28586 629338 28822 629574
rect 28266 589658 28502 589894
rect 28586 589658 28822 589894
rect 28266 589338 28502 589574
rect 28586 589338 28822 589574
rect 28266 549658 28502 549894
rect 28586 549658 28822 549894
rect 28266 549338 28502 549574
rect 28586 549338 28822 549574
rect 28266 509658 28502 509894
rect 28586 509658 28822 509894
rect 28266 509338 28502 509574
rect 28586 509338 28822 509574
rect 28266 469658 28502 469894
rect 28586 469658 28822 469894
rect 28266 469338 28502 469574
rect 28586 469338 28822 469574
rect 28266 429658 28502 429894
rect 28586 429658 28822 429894
rect 28266 429338 28502 429574
rect 28586 429338 28822 429574
rect 28266 389658 28502 389894
rect 28586 389658 28822 389894
rect 28266 389338 28502 389574
rect 28586 389338 28822 389574
rect 28266 349658 28502 349894
rect 28586 349658 28822 349894
rect 28266 349338 28502 349574
rect 28586 349338 28822 349574
rect 28266 309658 28502 309894
rect 28586 309658 28822 309894
rect 28266 309338 28502 309574
rect 28586 309338 28822 309574
rect 28266 269658 28502 269894
rect 28586 269658 28822 269894
rect 28266 269338 28502 269574
rect 28586 269338 28822 269574
rect 28266 229658 28502 229894
rect 28586 229658 28822 229894
rect 28266 229338 28502 229574
rect 28586 229338 28822 229574
rect 28266 189658 28502 189894
rect 28586 189658 28822 189894
rect 28266 189338 28502 189574
rect 28586 189338 28822 189574
rect 28266 149658 28502 149894
rect 28586 149658 28822 149894
rect 28266 149338 28502 149574
rect 28586 149338 28822 149574
rect 28266 109658 28502 109894
rect 28586 109658 28822 109894
rect 28266 109338 28502 109574
rect 28586 109338 28822 109574
rect 28266 69658 28502 69894
rect 28586 69658 28822 69894
rect 28266 69338 28502 69574
rect 28586 69338 28822 69574
rect 28266 29658 28502 29894
rect 28586 29658 28822 29894
rect 28266 29338 28502 29574
rect 28586 29338 28822 29574
rect 28266 -5382 28502 -5146
rect 28586 -5382 28822 -5146
rect 28266 -5702 28502 -5466
rect 28586 -5702 28822 -5466
rect 51986 710362 52222 710598
rect 52306 710362 52542 710598
rect 51986 710042 52222 710278
rect 52306 710042 52542 710278
rect 48266 708442 48502 708678
rect 48586 708442 48822 708678
rect 48266 708122 48502 708358
rect 48586 708122 48822 708358
rect 44546 706522 44782 706758
rect 44866 706522 45102 706758
rect 44546 706202 44782 706438
rect 44866 706202 45102 706438
rect 31986 673378 32222 673614
rect 32306 673378 32542 673614
rect 31986 673058 32222 673294
rect 32306 673058 32542 673294
rect 31986 633378 32222 633614
rect 32306 633378 32542 633614
rect 31986 633058 32222 633294
rect 32306 633058 32542 633294
rect 31986 593378 32222 593614
rect 32306 593378 32542 593614
rect 31986 593058 32222 593294
rect 32306 593058 32542 593294
rect 31986 553378 32222 553614
rect 32306 553378 32542 553614
rect 31986 553058 32222 553294
rect 32306 553058 32542 553294
rect 31986 513378 32222 513614
rect 32306 513378 32542 513614
rect 31986 513058 32222 513294
rect 32306 513058 32542 513294
rect 31986 473378 32222 473614
rect 32306 473378 32542 473614
rect 31986 473058 32222 473294
rect 32306 473058 32542 473294
rect 31986 433378 32222 433614
rect 32306 433378 32542 433614
rect 31986 433058 32222 433294
rect 32306 433058 32542 433294
rect 31986 393378 32222 393614
rect 32306 393378 32542 393614
rect 31986 393058 32222 393294
rect 32306 393058 32542 393294
rect 31986 353378 32222 353614
rect 32306 353378 32542 353614
rect 31986 353058 32222 353294
rect 32306 353058 32542 353294
rect 31986 313378 32222 313614
rect 32306 313378 32542 313614
rect 31986 313058 32222 313294
rect 32306 313058 32542 313294
rect 31986 273378 32222 273614
rect 32306 273378 32542 273614
rect 31986 273058 32222 273294
rect 32306 273058 32542 273294
rect 31986 233378 32222 233614
rect 32306 233378 32542 233614
rect 31986 233058 32222 233294
rect 32306 233058 32542 233294
rect 31986 193378 32222 193614
rect 32306 193378 32542 193614
rect 31986 193058 32222 193294
rect 32306 193058 32542 193294
rect 31986 153378 32222 153614
rect 32306 153378 32542 153614
rect 31986 153058 32222 153294
rect 32306 153058 32542 153294
rect 31986 113378 32222 113614
rect 32306 113378 32542 113614
rect 31986 113058 32222 113294
rect 32306 113058 32542 113294
rect 31986 73378 32222 73614
rect 32306 73378 32542 73614
rect 31986 73058 32222 73294
rect 32306 73058 32542 73294
rect 31986 33378 32222 33614
rect 32306 33378 32542 33614
rect 31986 33058 32222 33294
rect 32306 33058 32542 33294
rect 11986 -6342 12222 -6106
rect 12306 -6342 12542 -6106
rect 11986 -6662 12222 -6426
rect 12306 -6662 12542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 40826 704602 41062 704838
rect 41146 704602 41382 704838
rect 40826 704282 41062 704518
rect 41146 704282 41382 704518
rect 40826 682218 41062 682454
rect 41146 682218 41382 682454
rect 40826 681898 41062 682134
rect 41146 681898 41382 682134
rect 40826 642218 41062 642454
rect 41146 642218 41382 642454
rect 40826 641898 41062 642134
rect 41146 641898 41382 642134
rect 40826 602218 41062 602454
rect 41146 602218 41382 602454
rect 40826 601898 41062 602134
rect 41146 601898 41382 602134
rect 40826 562218 41062 562454
rect 41146 562218 41382 562454
rect 40826 561898 41062 562134
rect 41146 561898 41382 562134
rect 40826 522218 41062 522454
rect 41146 522218 41382 522454
rect 40826 521898 41062 522134
rect 41146 521898 41382 522134
rect 40826 482218 41062 482454
rect 41146 482218 41382 482454
rect 40826 481898 41062 482134
rect 41146 481898 41382 482134
rect 40826 442218 41062 442454
rect 41146 442218 41382 442454
rect 40826 441898 41062 442134
rect 41146 441898 41382 442134
rect 40826 402218 41062 402454
rect 41146 402218 41382 402454
rect 40826 401898 41062 402134
rect 41146 401898 41382 402134
rect 40826 362218 41062 362454
rect 41146 362218 41382 362454
rect 40826 361898 41062 362134
rect 41146 361898 41382 362134
rect 40826 322218 41062 322454
rect 41146 322218 41382 322454
rect 40826 321898 41062 322134
rect 41146 321898 41382 322134
rect 40826 282218 41062 282454
rect 41146 282218 41382 282454
rect 40826 281898 41062 282134
rect 41146 281898 41382 282134
rect 40826 242218 41062 242454
rect 41146 242218 41382 242454
rect 40826 241898 41062 242134
rect 41146 241898 41382 242134
rect 40826 202218 41062 202454
rect 41146 202218 41382 202454
rect 40826 201898 41062 202134
rect 41146 201898 41382 202134
rect 40826 162218 41062 162454
rect 41146 162218 41382 162454
rect 40826 161898 41062 162134
rect 41146 161898 41382 162134
rect 40826 122218 41062 122454
rect 41146 122218 41382 122454
rect 40826 121898 41062 122134
rect 41146 121898 41382 122134
rect 40826 82218 41062 82454
rect 41146 82218 41382 82454
rect 40826 81898 41062 82134
rect 41146 81898 41382 82134
rect 40826 42218 41062 42454
rect 41146 42218 41382 42454
rect 40826 41898 41062 42134
rect 41146 41898 41382 42134
rect 40826 2218 41062 2454
rect 41146 2218 41382 2454
rect 40826 1898 41062 2134
rect 41146 1898 41382 2134
rect 40826 -582 41062 -346
rect 41146 -582 41382 -346
rect 40826 -902 41062 -666
rect 41146 -902 41382 -666
rect 44546 685938 44782 686174
rect 44866 685938 45102 686174
rect 44546 685618 44782 685854
rect 44866 685618 45102 685854
rect 44546 645938 44782 646174
rect 44866 645938 45102 646174
rect 44546 645618 44782 645854
rect 44866 645618 45102 645854
rect 44546 605938 44782 606174
rect 44866 605938 45102 606174
rect 44546 605618 44782 605854
rect 44866 605618 45102 605854
rect 44546 565938 44782 566174
rect 44866 565938 45102 566174
rect 44546 565618 44782 565854
rect 44866 565618 45102 565854
rect 44546 525938 44782 526174
rect 44866 525938 45102 526174
rect 44546 525618 44782 525854
rect 44866 525618 45102 525854
rect 44546 485938 44782 486174
rect 44866 485938 45102 486174
rect 44546 485618 44782 485854
rect 44866 485618 45102 485854
rect 44546 445938 44782 446174
rect 44866 445938 45102 446174
rect 44546 445618 44782 445854
rect 44866 445618 45102 445854
rect 44546 405938 44782 406174
rect 44866 405938 45102 406174
rect 44546 405618 44782 405854
rect 44866 405618 45102 405854
rect 44546 365938 44782 366174
rect 44866 365938 45102 366174
rect 44546 365618 44782 365854
rect 44866 365618 45102 365854
rect 44546 325938 44782 326174
rect 44866 325938 45102 326174
rect 44546 325618 44782 325854
rect 44866 325618 45102 325854
rect 44546 285938 44782 286174
rect 44866 285938 45102 286174
rect 44546 285618 44782 285854
rect 44866 285618 45102 285854
rect 44546 245938 44782 246174
rect 44866 245938 45102 246174
rect 44546 245618 44782 245854
rect 44866 245618 45102 245854
rect 44546 205938 44782 206174
rect 44866 205938 45102 206174
rect 44546 205618 44782 205854
rect 44866 205618 45102 205854
rect 44546 165938 44782 166174
rect 44866 165938 45102 166174
rect 44546 165618 44782 165854
rect 44866 165618 45102 165854
rect 44546 125938 44782 126174
rect 44866 125938 45102 126174
rect 44546 125618 44782 125854
rect 44866 125618 45102 125854
rect 44546 85938 44782 86174
rect 44866 85938 45102 86174
rect 44546 85618 44782 85854
rect 44866 85618 45102 85854
rect 44546 45938 44782 46174
rect 44866 45938 45102 46174
rect 44546 45618 44782 45854
rect 44866 45618 45102 45854
rect 44546 5938 44782 6174
rect 44866 5938 45102 6174
rect 44546 5618 44782 5854
rect 44866 5618 45102 5854
rect 44546 -2502 44782 -2266
rect 44866 -2502 45102 -2266
rect 44546 -2822 44782 -2586
rect 44866 -2822 45102 -2586
rect 48266 689658 48502 689894
rect 48586 689658 48822 689894
rect 48266 689338 48502 689574
rect 48586 689338 48822 689574
rect 48266 649658 48502 649894
rect 48586 649658 48822 649894
rect 48266 649338 48502 649574
rect 48586 649338 48822 649574
rect 48266 609658 48502 609894
rect 48586 609658 48822 609894
rect 48266 609338 48502 609574
rect 48586 609338 48822 609574
rect 48266 569658 48502 569894
rect 48586 569658 48822 569894
rect 48266 569338 48502 569574
rect 48586 569338 48822 569574
rect 48266 529658 48502 529894
rect 48586 529658 48822 529894
rect 48266 529338 48502 529574
rect 48586 529338 48822 529574
rect 48266 489658 48502 489894
rect 48586 489658 48822 489894
rect 48266 489338 48502 489574
rect 48586 489338 48822 489574
rect 48266 449658 48502 449894
rect 48586 449658 48822 449894
rect 48266 449338 48502 449574
rect 48586 449338 48822 449574
rect 48266 409658 48502 409894
rect 48586 409658 48822 409894
rect 48266 409338 48502 409574
rect 48586 409338 48822 409574
rect 48266 369658 48502 369894
rect 48586 369658 48822 369894
rect 48266 369338 48502 369574
rect 48586 369338 48822 369574
rect 48266 329658 48502 329894
rect 48586 329658 48822 329894
rect 48266 329338 48502 329574
rect 48586 329338 48822 329574
rect 48266 289658 48502 289894
rect 48586 289658 48822 289894
rect 48266 289338 48502 289574
rect 48586 289338 48822 289574
rect 48266 249658 48502 249894
rect 48586 249658 48822 249894
rect 48266 249338 48502 249574
rect 48586 249338 48822 249574
rect 48266 209658 48502 209894
rect 48586 209658 48822 209894
rect 48266 209338 48502 209574
rect 48586 209338 48822 209574
rect 48266 169658 48502 169894
rect 48586 169658 48822 169894
rect 48266 169338 48502 169574
rect 48586 169338 48822 169574
rect 48266 129658 48502 129894
rect 48586 129658 48822 129894
rect 48266 129338 48502 129574
rect 48586 129338 48822 129574
rect 48266 89658 48502 89894
rect 48586 89658 48822 89894
rect 48266 89338 48502 89574
rect 48586 89338 48822 89574
rect 48266 49658 48502 49894
rect 48586 49658 48822 49894
rect 48266 49338 48502 49574
rect 48586 49338 48822 49574
rect 48266 9658 48502 9894
rect 48586 9658 48822 9894
rect 48266 9338 48502 9574
rect 48586 9338 48822 9574
rect 48266 -4422 48502 -4186
rect 48586 -4422 48822 -4186
rect 48266 -4742 48502 -4506
rect 48586 -4742 48822 -4506
rect 71986 711322 72222 711558
rect 72306 711322 72542 711558
rect 71986 711002 72222 711238
rect 72306 711002 72542 711238
rect 68266 709402 68502 709638
rect 68586 709402 68822 709638
rect 68266 709082 68502 709318
rect 68586 709082 68822 709318
rect 64546 707482 64782 707718
rect 64866 707482 65102 707718
rect 64546 707162 64782 707398
rect 64866 707162 65102 707398
rect 51986 693378 52222 693614
rect 52306 693378 52542 693614
rect 51986 693058 52222 693294
rect 52306 693058 52542 693294
rect 51986 653378 52222 653614
rect 52306 653378 52542 653614
rect 51986 653058 52222 653294
rect 52306 653058 52542 653294
rect 51986 613378 52222 613614
rect 52306 613378 52542 613614
rect 51986 613058 52222 613294
rect 52306 613058 52542 613294
rect 51986 573378 52222 573614
rect 52306 573378 52542 573614
rect 51986 573058 52222 573294
rect 52306 573058 52542 573294
rect 51986 533378 52222 533614
rect 52306 533378 52542 533614
rect 51986 533058 52222 533294
rect 52306 533058 52542 533294
rect 51986 493378 52222 493614
rect 52306 493378 52542 493614
rect 51986 493058 52222 493294
rect 52306 493058 52542 493294
rect 51986 453378 52222 453614
rect 52306 453378 52542 453614
rect 51986 453058 52222 453294
rect 52306 453058 52542 453294
rect 51986 413378 52222 413614
rect 52306 413378 52542 413614
rect 51986 413058 52222 413294
rect 52306 413058 52542 413294
rect 51986 373378 52222 373614
rect 52306 373378 52542 373614
rect 51986 373058 52222 373294
rect 52306 373058 52542 373294
rect 51986 333378 52222 333614
rect 52306 333378 52542 333614
rect 51986 333058 52222 333294
rect 52306 333058 52542 333294
rect 51986 293378 52222 293614
rect 52306 293378 52542 293614
rect 51986 293058 52222 293294
rect 52306 293058 52542 293294
rect 51986 253378 52222 253614
rect 52306 253378 52542 253614
rect 51986 253058 52222 253294
rect 52306 253058 52542 253294
rect 51986 213378 52222 213614
rect 52306 213378 52542 213614
rect 51986 213058 52222 213294
rect 52306 213058 52542 213294
rect 51986 173378 52222 173614
rect 52306 173378 52542 173614
rect 51986 173058 52222 173294
rect 52306 173058 52542 173294
rect 51986 133378 52222 133614
rect 52306 133378 52542 133614
rect 51986 133058 52222 133294
rect 52306 133058 52542 133294
rect 51986 93378 52222 93614
rect 52306 93378 52542 93614
rect 51986 93058 52222 93294
rect 52306 93058 52542 93294
rect 51986 53378 52222 53614
rect 52306 53378 52542 53614
rect 51986 53058 52222 53294
rect 52306 53058 52542 53294
rect 51986 13378 52222 13614
rect 52306 13378 52542 13614
rect 51986 13058 52222 13294
rect 52306 13058 52542 13294
rect 31986 -7302 32222 -7066
rect 32306 -7302 32542 -7066
rect 31986 -7622 32222 -7386
rect 32306 -7622 32542 -7386
rect 60826 705562 61062 705798
rect 61146 705562 61382 705798
rect 60826 705242 61062 705478
rect 61146 705242 61382 705478
rect 60826 662218 61062 662454
rect 61146 662218 61382 662454
rect 60826 661898 61062 662134
rect 61146 661898 61382 662134
rect 60826 622218 61062 622454
rect 61146 622218 61382 622454
rect 60826 621898 61062 622134
rect 61146 621898 61382 622134
rect 60826 582218 61062 582454
rect 61146 582218 61382 582454
rect 60826 581898 61062 582134
rect 61146 581898 61382 582134
rect 60826 542218 61062 542454
rect 61146 542218 61382 542454
rect 60826 541898 61062 542134
rect 61146 541898 61382 542134
rect 60826 502218 61062 502454
rect 61146 502218 61382 502454
rect 60826 501898 61062 502134
rect 61146 501898 61382 502134
rect 60826 462218 61062 462454
rect 61146 462218 61382 462454
rect 60826 461898 61062 462134
rect 61146 461898 61382 462134
rect 60826 422218 61062 422454
rect 61146 422218 61382 422454
rect 60826 421898 61062 422134
rect 61146 421898 61382 422134
rect 60826 382218 61062 382454
rect 61146 382218 61382 382454
rect 60826 381898 61062 382134
rect 61146 381898 61382 382134
rect 60826 342218 61062 342454
rect 61146 342218 61382 342454
rect 60826 341898 61062 342134
rect 61146 341898 61382 342134
rect 60826 302218 61062 302454
rect 61146 302218 61382 302454
rect 60826 301898 61062 302134
rect 61146 301898 61382 302134
rect 60826 262218 61062 262454
rect 61146 262218 61382 262454
rect 60826 261898 61062 262134
rect 61146 261898 61382 262134
rect 60826 222218 61062 222454
rect 61146 222218 61382 222454
rect 60826 221898 61062 222134
rect 61146 221898 61382 222134
rect 60826 182218 61062 182454
rect 61146 182218 61382 182454
rect 60826 181898 61062 182134
rect 61146 181898 61382 182134
rect 60826 142218 61062 142454
rect 61146 142218 61382 142454
rect 60826 141898 61062 142134
rect 61146 141898 61382 142134
rect 60826 102218 61062 102454
rect 61146 102218 61382 102454
rect 60826 101898 61062 102134
rect 61146 101898 61382 102134
rect 60826 62218 61062 62454
rect 61146 62218 61382 62454
rect 60826 61898 61062 62134
rect 61146 61898 61382 62134
rect 60826 22218 61062 22454
rect 61146 22218 61382 22454
rect 60826 21898 61062 22134
rect 61146 21898 61382 22134
rect 60826 -1542 61062 -1306
rect 61146 -1542 61382 -1306
rect 60826 -1862 61062 -1626
rect 61146 -1862 61382 -1626
rect 64546 665938 64782 666174
rect 64866 665938 65102 666174
rect 64546 665618 64782 665854
rect 64866 665618 65102 665854
rect 64546 625938 64782 626174
rect 64866 625938 65102 626174
rect 64546 625618 64782 625854
rect 64866 625618 65102 625854
rect 64546 585938 64782 586174
rect 64866 585938 65102 586174
rect 64546 585618 64782 585854
rect 64866 585618 65102 585854
rect 64546 545938 64782 546174
rect 64866 545938 65102 546174
rect 64546 545618 64782 545854
rect 64866 545618 65102 545854
rect 64546 505938 64782 506174
rect 64866 505938 65102 506174
rect 64546 505618 64782 505854
rect 64866 505618 65102 505854
rect 64546 465938 64782 466174
rect 64866 465938 65102 466174
rect 64546 465618 64782 465854
rect 64866 465618 65102 465854
rect 64546 425938 64782 426174
rect 64866 425938 65102 426174
rect 64546 425618 64782 425854
rect 64866 425618 65102 425854
rect 64546 385938 64782 386174
rect 64866 385938 65102 386174
rect 64546 385618 64782 385854
rect 64866 385618 65102 385854
rect 64546 345938 64782 346174
rect 64866 345938 65102 346174
rect 64546 345618 64782 345854
rect 64866 345618 65102 345854
rect 64546 305938 64782 306174
rect 64866 305938 65102 306174
rect 64546 305618 64782 305854
rect 64866 305618 65102 305854
rect 64546 265938 64782 266174
rect 64866 265938 65102 266174
rect 64546 265618 64782 265854
rect 64866 265618 65102 265854
rect 64546 225938 64782 226174
rect 64866 225938 65102 226174
rect 64546 225618 64782 225854
rect 64866 225618 65102 225854
rect 64546 185938 64782 186174
rect 64866 185938 65102 186174
rect 64546 185618 64782 185854
rect 64866 185618 65102 185854
rect 64546 145938 64782 146174
rect 64866 145938 65102 146174
rect 64546 145618 64782 145854
rect 64866 145618 65102 145854
rect 64546 105938 64782 106174
rect 64866 105938 65102 106174
rect 64546 105618 64782 105854
rect 64866 105618 65102 105854
rect 64546 65938 64782 66174
rect 64866 65938 65102 66174
rect 64546 65618 64782 65854
rect 64866 65618 65102 65854
rect 64546 25938 64782 26174
rect 64866 25938 65102 26174
rect 64546 25618 64782 25854
rect 64866 25618 65102 25854
rect 64546 -3462 64782 -3226
rect 64866 -3462 65102 -3226
rect 64546 -3782 64782 -3546
rect 64866 -3782 65102 -3546
rect 68266 669658 68502 669894
rect 68586 669658 68822 669894
rect 68266 669338 68502 669574
rect 68586 669338 68822 669574
rect 68266 629658 68502 629894
rect 68586 629658 68822 629894
rect 68266 629338 68502 629574
rect 68586 629338 68822 629574
rect 68266 589658 68502 589894
rect 68586 589658 68822 589894
rect 68266 589338 68502 589574
rect 68586 589338 68822 589574
rect 68266 549658 68502 549894
rect 68586 549658 68822 549894
rect 68266 549338 68502 549574
rect 68586 549338 68822 549574
rect 68266 509658 68502 509894
rect 68586 509658 68822 509894
rect 68266 509338 68502 509574
rect 68586 509338 68822 509574
rect 68266 469658 68502 469894
rect 68586 469658 68822 469894
rect 68266 469338 68502 469574
rect 68586 469338 68822 469574
rect 68266 429658 68502 429894
rect 68586 429658 68822 429894
rect 68266 429338 68502 429574
rect 68586 429338 68822 429574
rect 68266 389658 68502 389894
rect 68586 389658 68822 389894
rect 68266 389338 68502 389574
rect 68586 389338 68822 389574
rect 68266 349658 68502 349894
rect 68586 349658 68822 349894
rect 68266 349338 68502 349574
rect 68586 349338 68822 349574
rect 68266 309658 68502 309894
rect 68586 309658 68822 309894
rect 68266 309338 68502 309574
rect 68586 309338 68822 309574
rect 68266 269658 68502 269894
rect 68586 269658 68822 269894
rect 68266 269338 68502 269574
rect 68586 269338 68822 269574
rect 68266 229658 68502 229894
rect 68586 229658 68822 229894
rect 68266 229338 68502 229574
rect 68586 229338 68822 229574
rect 68266 189658 68502 189894
rect 68586 189658 68822 189894
rect 68266 189338 68502 189574
rect 68586 189338 68822 189574
rect 68266 149658 68502 149894
rect 68586 149658 68822 149894
rect 68266 149338 68502 149574
rect 68586 149338 68822 149574
rect 68266 109658 68502 109894
rect 68586 109658 68822 109894
rect 68266 109338 68502 109574
rect 68586 109338 68822 109574
rect 68266 69658 68502 69894
rect 68586 69658 68822 69894
rect 68266 69338 68502 69574
rect 68586 69338 68822 69574
rect 68266 29658 68502 29894
rect 68586 29658 68822 29894
rect 68266 29338 68502 29574
rect 68586 29338 68822 29574
rect 68266 -5382 68502 -5146
rect 68586 -5382 68822 -5146
rect 68266 -5702 68502 -5466
rect 68586 -5702 68822 -5466
rect 91986 710362 92222 710598
rect 92306 710362 92542 710598
rect 91986 710042 92222 710278
rect 92306 710042 92542 710278
rect 88266 708442 88502 708678
rect 88586 708442 88822 708678
rect 88266 708122 88502 708358
rect 88586 708122 88822 708358
rect 84546 706522 84782 706758
rect 84866 706522 85102 706758
rect 84546 706202 84782 706438
rect 84866 706202 85102 706438
rect 71986 673378 72222 673614
rect 72306 673378 72542 673614
rect 71986 673058 72222 673294
rect 72306 673058 72542 673294
rect 71986 633378 72222 633614
rect 72306 633378 72542 633614
rect 71986 633058 72222 633294
rect 72306 633058 72542 633294
rect 71986 593378 72222 593614
rect 72306 593378 72542 593614
rect 71986 593058 72222 593294
rect 72306 593058 72542 593294
rect 71986 553378 72222 553614
rect 72306 553378 72542 553614
rect 71986 553058 72222 553294
rect 72306 553058 72542 553294
rect 71986 513378 72222 513614
rect 72306 513378 72542 513614
rect 71986 513058 72222 513294
rect 72306 513058 72542 513294
rect 71986 473378 72222 473614
rect 72306 473378 72542 473614
rect 71986 473058 72222 473294
rect 72306 473058 72542 473294
rect 71986 433378 72222 433614
rect 72306 433378 72542 433614
rect 71986 433058 72222 433294
rect 72306 433058 72542 433294
rect 71986 393378 72222 393614
rect 72306 393378 72542 393614
rect 71986 393058 72222 393294
rect 72306 393058 72542 393294
rect 71986 353378 72222 353614
rect 72306 353378 72542 353614
rect 71986 353058 72222 353294
rect 72306 353058 72542 353294
rect 71986 313378 72222 313614
rect 72306 313378 72542 313614
rect 71986 313058 72222 313294
rect 72306 313058 72542 313294
rect 71986 273378 72222 273614
rect 72306 273378 72542 273614
rect 71986 273058 72222 273294
rect 72306 273058 72542 273294
rect 71986 233378 72222 233614
rect 72306 233378 72542 233614
rect 71986 233058 72222 233294
rect 72306 233058 72542 233294
rect 71986 193378 72222 193614
rect 72306 193378 72542 193614
rect 71986 193058 72222 193294
rect 72306 193058 72542 193294
rect 71986 153378 72222 153614
rect 72306 153378 72542 153614
rect 71986 153058 72222 153294
rect 72306 153058 72542 153294
rect 71986 113378 72222 113614
rect 72306 113378 72542 113614
rect 71986 113058 72222 113294
rect 72306 113058 72542 113294
rect 71986 73378 72222 73614
rect 72306 73378 72542 73614
rect 71986 73058 72222 73294
rect 72306 73058 72542 73294
rect 71986 33378 72222 33614
rect 72306 33378 72542 33614
rect 71986 33058 72222 33294
rect 72306 33058 72542 33294
rect 51986 -6342 52222 -6106
rect 52306 -6342 52542 -6106
rect 51986 -6662 52222 -6426
rect 52306 -6662 52542 -6426
rect 80826 704602 81062 704838
rect 81146 704602 81382 704838
rect 80826 704282 81062 704518
rect 81146 704282 81382 704518
rect 80826 682218 81062 682454
rect 81146 682218 81382 682454
rect 80826 681898 81062 682134
rect 81146 681898 81382 682134
rect 80826 642218 81062 642454
rect 81146 642218 81382 642454
rect 80826 641898 81062 642134
rect 81146 641898 81382 642134
rect 80826 602218 81062 602454
rect 81146 602218 81382 602454
rect 80826 601898 81062 602134
rect 81146 601898 81382 602134
rect 80826 562218 81062 562454
rect 81146 562218 81382 562454
rect 80826 561898 81062 562134
rect 81146 561898 81382 562134
rect 80826 522218 81062 522454
rect 81146 522218 81382 522454
rect 80826 521898 81062 522134
rect 81146 521898 81382 522134
rect 80826 482218 81062 482454
rect 81146 482218 81382 482454
rect 80826 481898 81062 482134
rect 81146 481898 81382 482134
rect 80826 442218 81062 442454
rect 81146 442218 81382 442454
rect 80826 441898 81062 442134
rect 81146 441898 81382 442134
rect 80826 402218 81062 402454
rect 81146 402218 81382 402454
rect 80826 401898 81062 402134
rect 81146 401898 81382 402134
rect 80826 362218 81062 362454
rect 81146 362218 81382 362454
rect 80826 361898 81062 362134
rect 81146 361898 81382 362134
rect 80826 322218 81062 322454
rect 81146 322218 81382 322454
rect 80826 321898 81062 322134
rect 81146 321898 81382 322134
rect 80826 282218 81062 282454
rect 81146 282218 81382 282454
rect 80826 281898 81062 282134
rect 81146 281898 81382 282134
rect 80826 242218 81062 242454
rect 81146 242218 81382 242454
rect 80826 241898 81062 242134
rect 81146 241898 81382 242134
rect 80826 202218 81062 202454
rect 81146 202218 81382 202454
rect 80826 201898 81062 202134
rect 81146 201898 81382 202134
rect 80826 162218 81062 162454
rect 81146 162218 81382 162454
rect 80826 161898 81062 162134
rect 81146 161898 81382 162134
rect 80826 122218 81062 122454
rect 81146 122218 81382 122454
rect 80826 121898 81062 122134
rect 81146 121898 81382 122134
rect 80826 82218 81062 82454
rect 81146 82218 81382 82454
rect 80826 81898 81062 82134
rect 81146 81898 81382 82134
rect 80826 42218 81062 42454
rect 81146 42218 81382 42454
rect 80826 41898 81062 42134
rect 81146 41898 81382 42134
rect 80826 2218 81062 2454
rect 81146 2218 81382 2454
rect 80826 1898 81062 2134
rect 81146 1898 81382 2134
rect 80826 -582 81062 -346
rect 81146 -582 81382 -346
rect 80826 -902 81062 -666
rect 81146 -902 81382 -666
rect 84546 685938 84782 686174
rect 84866 685938 85102 686174
rect 84546 685618 84782 685854
rect 84866 685618 85102 685854
rect 84546 645938 84782 646174
rect 84866 645938 85102 646174
rect 84546 645618 84782 645854
rect 84866 645618 85102 645854
rect 84546 605938 84782 606174
rect 84866 605938 85102 606174
rect 84546 605618 84782 605854
rect 84866 605618 85102 605854
rect 84546 565938 84782 566174
rect 84866 565938 85102 566174
rect 84546 565618 84782 565854
rect 84866 565618 85102 565854
rect 84546 525938 84782 526174
rect 84866 525938 85102 526174
rect 84546 525618 84782 525854
rect 84866 525618 85102 525854
rect 84546 485938 84782 486174
rect 84866 485938 85102 486174
rect 84546 485618 84782 485854
rect 84866 485618 85102 485854
rect 84546 445938 84782 446174
rect 84866 445938 85102 446174
rect 84546 445618 84782 445854
rect 84866 445618 85102 445854
rect 84546 405938 84782 406174
rect 84866 405938 85102 406174
rect 84546 405618 84782 405854
rect 84866 405618 85102 405854
rect 84546 365938 84782 366174
rect 84866 365938 85102 366174
rect 84546 365618 84782 365854
rect 84866 365618 85102 365854
rect 84546 325938 84782 326174
rect 84866 325938 85102 326174
rect 84546 325618 84782 325854
rect 84866 325618 85102 325854
rect 84546 285938 84782 286174
rect 84866 285938 85102 286174
rect 84546 285618 84782 285854
rect 84866 285618 85102 285854
rect 84546 245938 84782 246174
rect 84866 245938 85102 246174
rect 84546 245618 84782 245854
rect 84866 245618 85102 245854
rect 84546 205938 84782 206174
rect 84866 205938 85102 206174
rect 84546 205618 84782 205854
rect 84866 205618 85102 205854
rect 84546 165938 84782 166174
rect 84866 165938 85102 166174
rect 84546 165618 84782 165854
rect 84866 165618 85102 165854
rect 84546 125938 84782 126174
rect 84866 125938 85102 126174
rect 84546 125618 84782 125854
rect 84866 125618 85102 125854
rect 84546 85938 84782 86174
rect 84866 85938 85102 86174
rect 84546 85618 84782 85854
rect 84866 85618 85102 85854
rect 84546 45938 84782 46174
rect 84866 45938 85102 46174
rect 84546 45618 84782 45854
rect 84866 45618 85102 45854
rect 84546 5938 84782 6174
rect 84866 5938 85102 6174
rect 84546 5618 84782 5854
rect 84866 5618 85102 5854
rect 84546 -2502 84782 -2266
rect 84866 -2502 85102 -2266
rect 84546 -2822 84782 -2586
rect 84866 -2822 85102 -2586
rect 88266 689658 88502 689894
rect 88586 689658 88822 689894
rect 88266 689338 88502 689574
rect 88586 689338 88822 689574
rect 88266 649658 88502 649894
rect 88586 649658 88822 649894
rect 88266 649338 88502 649574
rect 88586 649338 88822 649574
rect 88266 609658 88502 609894
rect 88586 609658 88822 609894
rect 88266 609338 88502 609574
rect 88586 609338 88822 609574
rect 88266 569658 88502 569894
rect 88586 569658 88822 569894
rect 88266 569338 88502 569574
rect 88586 569338 88822 569574
rect 88266 529658 88502 529894
rect 88586 529658 88822 529894
rect 88266 529338 88502 529574
rect 88586 529338 88822 529574
rect 88266 489658 88502 489894
rect 88586 489658 88822 489894
rect 88266 489338 88502 489574
rect 88586 489338 88822 489574
rect 88266 449658 88502 449894
rect 88586 449658 88822 449894
rect 88266 449338 88502 449574
rect 88586 449338 88822 449574
rect 88266 409658 88502 409894
rect 88586 409658 88822 409894
rect 88266 409338 88502 409574
rect 88586 409338 88822 409574
rect 88266 369658 88502 369894
rect 88586 369658 88822 369894
rect 88266 369338 88502 369574
rect 88586 369338 88822 369574
rect 88266 329658 88502 329894
rect 88586 329658 88822 329894
rect 88266 329338 88502 329574
rect 88586 329338 88822 329574
rect 88266 289658 88502 289894
rect 88586 289658 88822 289894
rect 88266 289338 88502 289574
rect 88586 289338 88822 289574
rect 88266 249658 88502 249894
rect 88586 249658 88822 249894
rect 88266 249338 88502 249574
rect 88586 249338 88822 249574
rect 88266 209658 88502 209894
rect 88586 209658 88822 209894
rect 88266 209338 88502 209574
rect 88586 209338 88822 209574
rect 88266 169658 88502 169894
rect 88586 169658 88822 169894
rect 88266 169338 88502 169574
rect 88586 169338 88822 169574
rect 88266 129658 88502 129894
rect 88586 129658 88822 129894
rect 88266 129338 88502 129574
rect 88586 129338 88822 129574
rect 88266 89658 88502 89894
rect 88586 89658 88822 89894
rect 88266 89338 88502 89574
rect 88586 89338 88822 89574
rect 88266 49658 88502 49894
rect 88586 49658 88822 49894
rect 88266 49338 88502 49574
rect 88586 49338 88822 49574
rect 88266 9658 88502 9894
rect 88586 9658 88822 9894
rect 88266 9338 88502 9574
rect 88586 9338 88822 9574
rect 88266 -4422 88502 -4186
rect 88586 -4422 88822 -4186
rect 88266 -4742 88502 -4506
rect 88586 -4742 88822 -4506
rect 111986 711322 112222 711558
rect 112306 711322 112542 711558
rect 111986 711002 112222 711238
rect 112306 711002 112542 711238
rect 108266 709402 108502 709638
rect 108586 709402 108822 709638
rect 108266 709082 108502 709318
rect 108586 709082 108822 709318
rect 104546 707482 104782 707718
rect 104866 707482 105102 707718
rect 104546 707162 104782 707398
rect 104866 707162 105102 707398
rect 91986 693378 92222 693614
rect 92306 693378 92542 693614
rect 91986 693058 92222 693294
rect 92306 693058 92542 693294
rect 91986 653378 92222 653614
rect 92306 653378 92542 653614
rect 91986 653058 92222 653294
rect 92306 653058 92542 653294
rect 91986 613378 92222 613614
rect 92306 613378 92542 613614
rect 91986 613058 92222 613294
rect 92306 613058 92542 613294
rect 91986 573378 92222 573614
rect 92306 573378 92542 573614
rect 91986 573058 92222 573294
rect 92306 573058 92542 573294
rect 91986 533378 92222 533614
rect 92306 533378 92542 533614
rect 91986 533058 92222 533294
rect 92306 533058 92542 533294
rect 91986 493378 92222 493614
rect 92306 493378 92542 493614
rect 91986 493058 92222 493294
rect 92306 493058 92542 493294
rect 91986 453378 92222 453614
rect 92306 453378 92542 453614
rect 91986 453058 92222 453294
rect 92306 453058 92542 453294
rect 91986 413378 92222 413614
rect 92306 413378 92542 413614
rect 91986 413058 92222 413294
rect 92306 413058 92542 413294
rect 91986 373378 92222 373614
rect 92306 373378 92542 373614
rect 91986 373058 92222 373294
rect 92306 373058 92542 373294
rect 91986 333378 92222 333614
rect 92306 333378 92542 333614
rect 91986 333058 92222 333294
rect 92306 333058 92542 333294
rect 91986 293378 92222 293614
rect 92306 293378 92542 293614
rect 91986 293058 92222 293294
rect 92306 293058 92542 293294
rect 91986 253378 92222 253614
rect 92306 253378 92542 253614
rect 91986 253058 92222 253294
rect 92306 253058 92542 253294
rect 91986 213378 92222 213614
rect 92306 213378 92542 213614
rect 91986 213058 92222 213294
rect 92306 213058 92542 213294
rect 91986 173378 92222 173614
rect 92306 173378 92542 173614
rect 91986 173058 92222 173294
rect 92306 173058 92542 173294
rect 91986 133378 92222 133614
rect 92306 133378 92542 133614
rect 91986 133058 92222 133294
rect 92306 133058 92542 133294
rect 91986 93378 92222 93614
rect 92306 93378 92542 93614
rect 91986 93058 92222 93294
rect 92306 93058 92542 93294
rect 91986 53378 92222 53614
rect 92306 53378 92542 53614
rect 91986 53058 92222 53294
rect 92306 53058 92542 53294
rect 91986 13378 92222 13614
rect 92306 13378 92542 13614
rect 91986 13058 92222 13294
rect 92306 13058 92542 13294
rect 71986 -7302 72222 -7066
rect 72306 -7302 72542 -7066
rect 71986 -7622 72222 -7386
rect 72306 -7622 72542 -7386
rect 100826 705562 101062 705798
rect 101146 705562 101382 705798
rect 100826 705242 101062 705478
rect 101146 705242 101382 705478
rect 100826 662218 101062 662454
rect 101146 662218 101382 662454
rect 100826 661898 101062 662134
rect 101146 661898 101382 662134
rect 100826 622218 101062 622454
rect 101146 622218 101382 622454
rect 100826 621898 101062 622134
rect 101146 621898 101382 622134
rect 100826 582218 101062 582454
rect 101146 582218 101382 582454
rect 100826 581898 101062 582134
rect 101146 581898 101382 582134
rect 100826 542218 101062 542454
rect 101146 542218 101382 542454
rect 100826 541898 101062 542134
rect 101146 541898 101382 542134
rect 100826 502218 101062 502454
rect 101146 502218 101382 502454
rect 100826 501898 101062 502134
rect 101146 501898 101382 502134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 422218 101062 422454
rect 101146 422218 101382 422454
rect 100826 421898 101062 422134
rect 101146 421898 101382 422134
rect 100826 382218 101062 382454
rect 101146 382218 101382 382454
rect 100826 381898 101062 382134
rect 101146 381898 101382 382134
rect 100826 342218 101062 342454
rect 101146 342218 101382 342454
rect 100826 341898 101062 342134
rect 101146 341898 101382 342134
rect 100826 302218 101062 302454
rect 101146 302218 101382 302454
rect 100826 301898 101062 302134
rect 101146 301898 101382 302134
rect 100826 262218 101062 262454
rect 101146 262218 101382 262454
rect 100826 261898 101062 262134
rect 101146 261898 101382 262134
rect 100826 222218 101062 222454
rect 101146 222218 101382 222454
rect 100826 221898 101062 222134
rect 101146 221898 101382 222134
rect 100826 182218 101062 182454
rect 101146 182218 101382 182454
rect 100826 181898 101062 182134
rect 101146 181898 101382 182134
rect 100826 142218 101062 142454
rect 101146 142218 101382 142454
rect 100826 141898 101062 142134
rect 101146 141898 101382 142134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 62218 101062 62454
rect 101146 62218 101382 62454
rect 100826 61898 101062 62134
rect 101146 61898 101382 62134
rect 100826 22218 101062 22454
rect 101146 22218 101382 22454
rect 100826 21898 101062 22134
rect 101146 21898 101382 22134
rect 100826 -1542 101062 -1306
rect 101146 -1542 101382 -1306
rect 100826 -1862 101062 -1626
rect 101146 -1862 101382 -1626
rect 104546 665938 104782 666174
rect 104866 665938 105102 666174
rect 104546 665618 104782 665854
rect 104866 665618 105102 665854
rect 104546 625938 104782 626174
rect 104866 625938 105102 626174
rect 104546 625618 104782 625854
rect 104866 625618 105102 625854
rect 104546 585938 104782 586174
rect 104866 585938 105102 586174
rect 104546 585618 104782 585854
rect 104866 585618 105102 585854
rect 104546 545938 104782 546174
rect 104866 545938 105102 546174
rect 104546 545618 104782 545854
rect 104866 545618 105102 545854
rect 104546 505938 104782 506174
rect 104866 505938 105102 506174
rect 104546 505618 104782 505854
rect 104866 505618 105102 505854
rect 104546 465938 104782 466174
rect 104866 465938 105102 466174
rect 104546 465618 104782 465854
rect 104866 465618 105102 465854
rect 104546 425938 104782 426174
rect 104866 425938 105102 426174
rect 104546 425618 104782 425854
rect 104866 425618 105102 425854
rect 104546 385938 104782 386174
rect 104866 385938 105102 386174
rect 104546 385618 104782 385854
rect 104866 385618 105102 385854
rect 104546 345938 104782 346174
rect 104866 345938 105102 346174
rect 104546 345618 104782 345854
rect 104866 345618 105102 345854
rect 104546 305938 104782 306174
rect 104866 305938 105102 306174
rect 104546 305618 104782 305854
rect 104866 305618 105102 305854
rect 104546 265938 104782 266174
rect 104866 265938 105102 266174
rect 104546 265618 104782 265854
rect 104866 265618 105102 265854
rect 104546 225938 104782 226174
rect 104866 225938 105102 226174
rect 104546 225618 104782 225854
rect 104866 225618 105102 225854
rect 104546 185938 104782 186174
rect 104866 185938 105102 186174
rect 104546 185618 104782 185854
rect 104866 185618 105102 185854
rect 104546 145938 104782 146174
rect 104866 145938 105102 146174
rect 104546 145618 104782 145854
rect 104866 145618 105102 145854
rect 104546 105938 104782 106174
rect 104866 105938 105102 106174
rect 104546 105618 104782 105854
rect 104866 105618 105102 105854
rect 104546 65938 104782 66174
rect 104866 65938 105102 66174
rect 104546 65618 104782 65854
rect 104866 65618 105102 65854
rect 104546 25938 104782 26174
rect 104866 25938 105102 26174
rect 104546 25618 104782 25854
rect 104866 25618 105102 25854
rect 104546 -3462 104782 -3226
rect 104866 -3462 105102 -3226
rect 104546 -3782 104782 -3546
rect 104866 -3782 105102 -3546
rect 108266 669658 108502 669894
rect 108586 669658 108822 669894
rect 108266 669338 108502 669574
rect 108586 669338 108822 669574
rect 108266 629658 108502 629894
rect 108586 629658 108822 629894
rect 108266 629338 108502 629574
rect 108586 629338 108822 629574
rect 108266 589658 108502 589894
rect 108586 589658 108822 589894
rect 108266 589338 108502 589574
rect 108586 589338 108822 589574
rect 108266 549658 108502 549894
rect 108586 549658 108822 549894
rect 108266 549338 108502 549574
rect 108586 549338 108822 549574
rect 108266 509658 108502 509894
rect 108586 509658 108822 509894
rect 108266 509338 108502 509574
rect 108586 509338 108822 509574
rect 108266 469658 108502 469894
rect 108586 469658 108822 469894
rect 108266 469338 108502 469574
rect 108586 469338 108822 469574
rect 108266 429658 108502 429894
rect 108586 429658 108822 429894
rect 108266 429338 108502 429574
rect 108586 429338 108822 429574
rect 108266 389658 108502 389894
rect 108586 389658 108822 389894
rect 108266 389338 108502 389574
rect 108586 389338 108822 389574
rect 108266 349658 108502 349894
rect 108586 349658 108822 349894
rect 108266 349338 108502 349574
rect 108586 349338 108822 349574
rect 108266 309658 108502 309894
rect 108586 309658 108822 309894
rect 108266 309338 108502 309574
rect 108586 309338 108822 309574
rect 108266 269658 108502 269894
rect 108586 269658 108822 269894
rect 108266 269338 108502 269574
rect 108586 269338 108822 269574
rect 108266 229658 108502 229894
rect 108586 229658 108822 229894
rect 108266 229338 108502 229574
rect 108586 229338 108822 229574
rect 108266 189658 108502 189894
rect 108586 189658 108822 189894
rect 108266 189338 108502 189574
rect 108586 189338 108822 189574
rect 108266 149658 108502 149894
rect 108586 149658 108822 149894
rect 108266 149338 108502 149574
rect 108586 149338 108822 149574
rect 108266 109658 108502 109894
rect 108586 109658 108822 109894
rect 108266 109338 108502 109574
rect 108586 109338 108822 109574
rect 108266 69658 108502 69894
rect 108586 69658 108822 69894
rect 108266 69338 108502 69574
rect 108586 69338 108822 69574
rect 108266 29658 108502 29894
rect 108586 29658 108822 29894
rect 108266 29338 108502 29574
rect 108586 29338 108822 29574
rect 108266 -5382 108502 -5146
rect 108586 -5382 108822 -5146
rect 108266 -5702 108502 -5466
rect 108586 -5702 108822 -5466
rect 131986 710362 132222 710598
rect 132306 710362 132542 710598
rect 131986 710042 132222 710278
rect 132306 710042 132542 710278
rect 128266 708442 128502 708678
rect 128586 708442 128822 708678
rect 128266 708122 128502 708358
rect 128586 708122 128822 708358
rect 124546 706522 124782 706758
rect 124866 706522 125102 706758
rect 124546 706202 124782 706438
rect 124866 706202 125102 706438
rect 111986 673378 112222 673614
rect 112306 673378 112542 673614
rect 111986 673058 112222 673294
rect 112306 673058 112542 673294
rect 111986 633378 112222 633614
rect 112306 633378 112542 633614
rect 111986 633058 112222 633294
rect 112306 633058 112542 633294
rect 111986 593378 112222 593614
rect 112306 593378 112542 593614
rect 111986 593058 112222 593294
rect 112306 593058 112542 593294
rect 111986 553378 112222 553614
rect 112306 553378 112542 553614
rect 111986 553058 112222 553294
rect 112306 553058 112542 553294
rect 111986 513378 112222 513614
rect 112306 513378 112542 513614
rect 111986 513058 112222 513294
rect 112306 513058 112542 513294
rect 111986 473378 112222 473614
rect 112306 473378 112542 473614
rect 111986 473058 112222 473294
rect 112306 473058 112542 473294
rect 111986 433378 112222 433614
rect 112306 433378 112542 433614
rect 111986 433058 112222 433294
rect 112306 433058 112542 433294
rect 111986 393378 112222 393614
rect 112306 393378 112542 393614
rect 111986 393058 112222 393294
rect 112306 393058 112542 393294
rect 111986 353378 112222 353614
rect 112306 353378 112542 353614
rect 111986 353058 112222 353294
rect 112306 353058 112542 353294
rect 111986 313378 112222 313614
rect 112306 313378 112542 313614
rect 111986 313058 112222 313294
rect 112306 313058 112542 313294
rect 111986 273378 112222 273614
rect 112306 273378 112542 273614
rect 111986 273058 112222 273294
rect 112306 273058 112542 273294
rect 111986 233378 112222 233614
rect 112306 233378 112542 233614
rect 111986 233058 112222 233294
rect 112306 233058 112542 233294
rect 111986 193378 112222 193614
rect 112306 193378 112542 193614
rect 111986 193058 112222 193294
rect 112306 193058 112542 193294
rect 111986 153378 112222 153614
rect 112306 153378 112542 153614
rect 111986 153058 112222 153294
rect 112306 153058 112542 153294
rect 111986 113378 112222 113614
rect 112306 113378 112542 113614
rect 111986 113058 112222 113294
rect 112306 113058 112542 113294
rect 111986 73378 112222 73614
rect 112306 73378 112542 73614
rect 111986 73058 112222 73294
rect 112306 73058 112542 73294
rect 111986 33378 112222 33614
rect 112306 33378 112542 33614
rect 111986 33058 112222 33294
rect 112306 33058 112542 33294
rect 91986 -6342 92222 -6106
rect 92306 -6342 92542 -6106
rect 91986 -6662 92222 -6426
rect 92306 -6662 92542 -6426
rect 120826 704602 121062 704838
rect 121146 704602 121382 704838
rect 120826 704282 121062 704518
rect 121146 704282 121382 704518
rect 120826 682218 121062 682454
rect 121146 682218 121382 682454
rect 120826 681898 121062 682134
rect 121146 681898 121382 682134
rect 120826 642218 121062 642454
rect 121146 642218 121382 642454
rect 120826 641898 121062 642134
rect 121146 641898 121382 642134
rect 120826 602218 121062 602454
rect 121146 602218 121382 602454
rect 120826 601898 121062 602134
rect 121146 601898 121382 602134
rect 120826 562218 121062 562454
rect 121146 562218 121382 562454
rect 120826 561898 121062 562134
rect 121146 561898 121382 562134
rect 120826 522218 121062 522454
rect 121146 522218 121382 522454
rect 120826 521898 121062 522134
rect 121146 521898 121382 522134
rect 120826 482218 121062 482454
rect 121146 482218 121382 482454
rect 120826 481898 121062 482134
rect 121146 481898 121382 482134
rect 120826 442218 121062 442454
rect 121146 442218 121382 442454
rect 120826 441898 121062 442134
rect 121146 441898 121382 442134
rect 120826 402218 121062 402454
rect 121146 402218 121382 402454
rect 120826 401898 121062 402134
rect 121146 401898 121382 402134
rect 120826 362218 121062 362454
rect 121146 362218 121382 362454
rect 120826 361898 121062 362134
rect 121146 361898 121382 362134
rect 120826 322218 121062 322454
rect 121146 322218 121382 322454
rect 120826 321898 121062 322134
rect 121146 321898 121382 322134
rect 120826 282218 121062 282454
rect 121146 282218 121382 282454
rect 120826 281898 121062 282134
rect 121146 281898 121382 282134
rect 120826 242218 121062 242454
rect 121146 242218 121382 242454
rect 120826 241898 121062 242134
rect 121146 241898 121382 242134
rect 120826 202218 121062 202454
rect 121146 202218 121382 202454
rect 120826 201898 121062 202134
rect 121146 201898 121382 202134
rect 120826 162218 121062 162454
rect 121146 162218 121382 162454
rect 120826 161898 121062 162134
rect 121146 161898 121382 162134
rect 120826 122218 121062 122454
rect 121146 122218 121382 122454
rect 120826 121898 121062 122134
rect 121146 121898 121382 122134
rect 120826 82218 121062 82454
rect 121146 82218 121382 82454
rect 120826 81898 121062 82134
rect 121146 81898 121382 82134
rect 120826 42218 121062 42454
rect 121146 42218 121382 42454
rect 120826 41898 121062 42134
rect 121146 41898 121382 42134
rect 120826 2218 121062 2454
rect 121146 2218 121382 2454
rect 120826 1898 121062 2134
rect 121146 1898 121382 2134
rect 120826 -582 121062 -346
rect 121146 -582 121382 -346
rect 120826 -902 121062 -666
rect 121146 -902 121382 -666
rect 124546 685938 124782 686174
rect 124866 685938 125102 686174
rect 124546 685618 124782 685854
rect 124866 685618 125102 685854
rect 124546 645938 124782 646174
rect 124866 645938 125102 646174
rect 124546 645618 124782 645854
rect 124866 645618 125102 645854
rect 124546 605938 124782 606174
rect 124866 605938 125102 606174
rect 124546 605618 124782 605854
rect 124866 605618 125102 605854
rect 124546 565938 124782 566174
rect 124866 565938 125102 566174
rect 124546 565618 124782 565854
rect 124866 565618 125102 565854
rect 124546 525938 124782 526174
rect 124866 525938 125102 526174
rect 124546 525618 124782 525854
rect 124866 525618 125102 525854
rect 124546 485938 124782 486174
rect 124866 485938 125102 486174
rect 124546 485618 124782 485854
rect 124866 485618 125102 485854
rect 124546 445938 124782 446174
rect 124866 445938 125102 446174
rect 124546 445618 124782 445854
rect 124866 445618 125102 445854
rect 124546 405938 124782 406174
rect 124866 405938 125102 406174
rect 124546 405618 124782 405854
rect 124866 405618 125102 405854
rect 124546 365938 124782 366174
rect 124866 365938 125102 366174
rect 124546 365618 124782 365854
rect 124866 365618 125102 365854
rect 124546 325938 124782 326174
rect 124866 325938 125102 326174
rect 124546 325618 124782 325854
rect 124866 325618 125102 325854
rect 124546 285938 124782 286174
rect 124866 285938 125102 286174
rect 124546 285618 124782 285854
rect 124866 285618 125102 285854
rect 124546 245938 124782 246174
rect 124866 245938 125102 246174
rect 124546 245618 124782 245854
rect 124866 245618 125102 245854
rect 124546 205938 124782 206174
rect 124866 205938 125102 206174
rect 124546 205618 124782 205854
rect 124866 205618 125102 205854
rect 124546 165938 124782 166174
rect 124866 165938 125102 166174
rect 124546 165618 124782 165854
rect 124866 165618 125102 165854
rect 124546 125938 124782 126174
rect 124866 125938 125102 126174
rect 124546 125618 124782 125854
rect 124866 125618 125102 125854
rect 124546 85938 124782 86174
rect 124866 85938 125102 86174
rect 124546 85618 124782 85854
rect 124866 85618 125102 85854
rect 124546 45938 124782 46174
rect 124866 45938 125102 46174
rect 124546 45618 124782 45854
rect 124866 45618 125102 45854
rect 124546 5938 124782 6174
rect 124866 5938 125102 6174
rect 124546 5618 124782 5854
rect 124866 5618 125102 5854
rect 124546 -2502 124782 -2266
rect 124866 -2502 125102 -2266
rect 124546 -2822 124782 -2586
rect 124866 -2822 125102 -2586
rect 128266 689658 128502 689894
rect 128586 689658 128822 689894
rect 128266 689338 128502 689574
rect 128586 689338 128822 689574
rect 128266 649658 128502 649894
rect 128586 649658 128822 649894
rect 128266 649338 128502 649574
rect 128586 649338 128822 649574
rect 128266 609658 128502 609894
rect 128586 609658 128822 609894
rect 128266 609338 128502 609574
rect 128586 609338 128822 609574
rect 128266 569658 128502 569894
rect 128586 569658 128822 569894
rect 128266 569338 128502 569574
rect 128586 569338 128822 569574
rect 128266 529658 128502 529894
rect 128586 529658 128822 529894
rect 128266 529338 128502 529574
rect 128586 529338 128822 529574
rect 128266 489658 128502 489894
rect 128586 489658 128822 489894
rect 128266 489338 128502 489574
rect 128586 489338 128822 489574
rect 128266 449658 128502 449894
rect 128586 449658 128822 449894
rect 128266 449338 128502 449574
rect 128586 449338 128822 449574
rect 128266 409658 128502 409894
rect 128586 409658 128822 409894
rect 128266 409338 128502 409574
rect 128586 409338 128822 409574
rect 128266 369658 128502 369894
rect 128586 369658 128822 369894
rect 128266 369338 128502 369574
rect 128586 369338 128822 369574
rect 128266 329658 128502 329894
rect 128586 329658 128822 329894
rect 128266 329338 128502 329574
rect 128586 329338 128822 329574
rect 128266 289658 128502 289894
rect 128586 289658 128822 289894
rect 128266 289338 128502 289574
rect 128586 289338 128822 289574
rect 128266 249658 128502 249894
rect 128586 249658 128822 249894
rect 128266 249338 128502 249574
rect 128586 249338 128822 249574
rect 128266 209658 128502 209894
rect 128586 209658 128822 209894
rect 128266 209338 128502 209574
rect 128586 209338 128822 209574
rect 128266 169658 128502 169894
rect 128586 169658 128822 169894
rect 128266 169338 128502 169574
rect 128586 169338 128822 169574
rect 128266 129658 128502 129894
rect 128586 129658 128822 129894
rect 128266 129338 128502 129574
rect 128586 129338 128822 129574
rect 128266 89658 128502 89894
rect 128586 89658 128822 89894
rect 128266 89338 128502 89574
rect 128586 89338 128822 89574
rect 128266 49658 128502 49894
rect 128586 49658 128822 49894
rect 128266 49338 128502 49574
rect 128586 49338 128822 49574
rect 128266 9658 128502 9894
rect 128586 9658 128822 9894
rect 128266 9338 128502 9574
rect 128586 9338 128822 9574
rect 128266 -4422 128502 -4186
rect 128586 -4422 128822 -4186
rect 128266 -4742 128502 -4506
rect 128586 -4742 128822 -4506
rect 151986 711322 152222 711558
rect 152306 711322 152542 711558
rect 151986 711002 152222 711238
rect 152306 711002 152542 711238
rect 148266 709402 148502 709638
rect 148586 709402 148822 709638
rect 148266 709082 148502 709318
rect 148586 709082 148822 709318
rect 144546 707482 144782 707718
rect 144866 707482 145102 707718
rect 144546 707162 144782 707398
rect 144866 707162 145102 707398
rect 131986 693378 132222 693614
rect 132306 693378 132542 693614
rect 131986 693058 132222 693294
rect 132306 693058 132542 693294
rect 131986 653378 132222 653614
rect 132306 653378 132542 653614
rect 131986 653058 132222 653294
rect 132306 653058 132542 653294
rect 131986 613378 132222 613614
rect 132306 613378 132542 613614
rect 131986 613058 132222 613294
rect 132306 613058 132542 613294
rect 131986 573378 132222 573614
rect 132306 573378 132542 573614
rect 131986 573058 132222 573294
rect 132306 573058 132542 573294
rect 131986 533378 132222 533614
rect 132306 533378 132542 533614
rect 131986 533058 132222 533294
rect 132306 533058 132542 533294
rect 131986 493378 132222 493614
rect 132306 493378 132542 493614
rect 131986 493058 132222 493294
rect 132306 493058 132542 493294
rect 131986 453378 132222 453614
rect 132306 453378 132542 453614
rect 131986 453058 132222 453294
rect 132306 453058 132542 453294
rect 131986 413378 132222 413614
rect 132306 413378 132542 413614
rect 131986 413058 132222 413294
rect 132306 413058 132542 413294
rect 131986 373378 132222 373614
rect 132306 373378 132542 373614
rect 131986 373058 132222 373294
rect 132306 373058 132542 373294
rect 131986 333378 132222 333614
rect 132306 333378 132542 333614
rect 131986 333058 132222 333294
rect 132306 333058 132542 333294
rect 140826 705562 141062 705798
rect 141146 705562 141382 705798
rect 140826 705242 141062 705478
rect 141146 705242 141382 705478
rect 140826 662218 141062 662454
rect 141146 662218 141382 662454
rect 140826 661898 141062 662134
rect 141146 661898 141382 662134
rect 140826 622218 141062 622454
rect 141146 622218 141382 622454
rect 140826 621898 141062 622134
rect 141146 621898 141382 622134
rect 140826 582218 141062 582454
rect 141146 582218 141382 582454
rect 140826 581898 141062 582134
rect 141146 581898 141382 582134
rect 140826 542218 141062 542454
rect 141146 542218 141382 542454
rect 140826 541898 141062 542134
rect 141146 541898 141382 542134
rect 140826 502218 141062 502454
rect 141146 502218 141382 502454
rect 140826 501898 141062 502134
rect 141146 501898 141382 502134
rect 140826 462218 141062 462454
rect 141146 462218 141382 462454
rect 140826 461898 141062 462134
rect 141146 461898 141382 462134
rect 140826 422218 141062 422454
rect 141146 422218 141382 422454
rect 140826 421898 141062 422134
rect 141146 421898 141382 422134
rect 140826 382218 141062 382454
rect 141146 382218 141382 382454
rect 140826 381898 141062 382134
rect 141146 381898 141382 382134
rect 140826 342218 141062 342454
rect 141146 342218 141382 342454
rect 140826 341898 141062 342134
rect 141146 341898 141382 342134
rect 131986 293378 132222 293614
rect 132306 293378 132542 293614
rect 131986 293058 132222 293294
rect 132306 293058 132542 293294
rect 131986 253378 132222 253614
rect 132306 253378 132542 253614
rect 131986 253058 132222 253294
rect 132306 253058 132542 253294
rect 131986 213378 132222 213614
rect 132306 213378 132542 213614
rect 131986 213058 132222 213294
rect 132306 213058 132542 213294
rect 131986 173378 132222 173614
rect 132306 173378 132542 173614
rect 131986 173058 132222 173294
rect 132306 173058 132542 173294
rect 131986 133378 132222 133614
rect 132306 133378 132542 133614
rect 131986 133058 132222 133294
rect 132306 133058 132542 133294
rect 131986 93378 132222 93614
rect 132306 93378 132542 93614
rect 131986 93058 132222 93294
rect 132306 93058 132542 93294
rect 131986 53378 132222 53614
rect 132306 53378 132542 53614
rect 131986 53058 132222 53294
rect 132306 53058 132542 53294
rect 131986 13378 132222 13614
rect 132306 13378 132542 13614
rect 131986 13058 132222 13294
rect 132306 13058 132542 13294
rect 111986 -7302 112222 -7066
rect 112306 -7302 112542 -7066
rect 111986 -7622 112222 -7386
rect 112306 -7622 112542 -7386
rect 140826 302218 141382 302454
rect 140826 301898 141382 302134
rect 140826 262218 141382 262454
rect 140826 261898 141382 262134
rect 140826 222218 141382 222454
rect 140826 221898 141382 222134
rect 140826 182218 141382 182454
rect 140826 181898 141382 182134
rect 140826 142218 141382 142454
rect 140826 141898 141382 142134
rect 140826 102218 141062 102454
rect 141146 102218 141382 102454
rect 140826 101898 141062 102134
rect 141146 101898 141382 102134
rect 140826 62218 141062 62454
rect 141146 62218 141382 62454
rect 140826 61898 141062 62134
rect 141146 61898 141382 62134
rect 140826 22218 141062 22454
rect 141146 22218 141382 22454
rect 140826 21898 141062 22134
rect 141146 21898 141382 22134
rect 140826 -1542 141062 -1306
rect 141146 -1542 141382 -1306
rect 140826 -1862 141062 -1626
rect 141146 -1862 141382 -1626
rect 144546 665938 144782 666174
rect 144866 665938 145102 666174
rect 144546 665618 144782 665854
rect 144866 665618 145102 665854
rect 144546 625938 144782 626174
rect 144866 625938 145102 626174
rect 144546 625618 144782 625854
rect 144866 625618 145102 625854
rect 144546 585938 144782 586174
rect 144866 585938 145102 586174
rect 144546 585618 144782 585854
rect 144866 585618 145102 585854
rect 144546 545938 144782 546174
rect 144866 545938 145102 546174
rect 144546 545618 144782 545854
rect 144866 545618 145102 545854
rect 144546 505938 144782 506174
rect 144866 505938 145102 506174
rect 144546 505618 144782 505854
rect 144866 505618 145102 505854
rect 144546 465938 144782 466174
rect 144866 465938 145102 466174
rect 144546 465618 144782 465854
rect 144866 465618 145102 465854
rect 144546 425938 144782 426174
rect 144866 425938 145102 426174
rect 144546 425618 144782 425854
rect 144866 425618 145102 425854
rect 144546 385938 144782 386174
rect 144866 385938 145102 386174
rect 144546 385618 144782 385854
rect 144866 385618 145102 385854
rect 144546 345938 144782 346174
rect 144866 345938 145102 346174
rect 144546 345618 144782 345854
rect 144866 345618 145102 345854
rect 144546 305938 144782 306174
rect 144866 305938 145102 306174
rect 144546 305618 144782 305854
rect 144866 305618 145102 305854
rect 144546 265938 144782 266174
rect 144866 265938 145102 266174
rect 144546 265618 144782 265854
rect 144866 265618 145102 265854
rect 144546 225938 144782 226174
rect 144866 225938 145102 226174
rect 144546 225618 144782 225854
rect 144866 225618 145102 225854
rect 144546 185938 144782 186174
rect 144866 185938 145102 186174
rect 144546 185618 144782 185854
rect 144866 185618 145102 185854
rect 144546 145938 144782 146174
rect 144866 145938 145102 146174
rect 144546 145618 144782 145854
rect 144866 145618 145102 145854
rect 144546 105938 144782 106174
rect 144866 105938 145102 106174
rect 144546 105618 144782 105854
rect 144866 105618 145102 105854
rect 144546 65938 144782 66174
rect 144866 65938 145102 66174
rect 144546 65618 144782 65854
rect 144866 65618 145102 65854
rect 144546 25938 144782 26174
rect 144866 25938 145102 26174
rect 144546 25618 144782 25854
rect 144866 25618 145102 25854
rect 144546 -3462 144782 -3226
rect 144866 -3462 145102 -3226
rect 144546 -3782 144782 -3546
rect 144866 -3782 145102 -3546
rect 148266 669658 148502 669894
rect 148586 669658 148822 669894
rect 148266 669338 148502 669574
rect 148586 669338 148822 669574
rect 148266 629658 148502 629894
rect 148586 629658 148822 629894
rect 148266 629338 148502 629574
rect 148586 629338 148822 629574
rect 148266 589658 148502 589894
rect 148586 589658 148822 589894
rect 148266 589338 148502 589574
rect 148586 589338 148822 589574
rect 148266 549658 148502 549894
rect 148586 549658 148822 549894
rect 148266 549338 148502 549574
rect 148586 549338 148822 549574
rect 148266 509658 148502 509894
rect 148586 509658 148822 509894
rect 148266 509338 148502 509574
rect 148586 509338 148822 509574
rect 148266 469658 148502 469894
rect 148586 469658 148822 469894
rect 148266 469338 148502 469574
rect 148586 469338 148822 469574
rect 148266 429658 148502 429894
rect 148586 429658 148822 429894
rect 148266 429338 148502 429574
rect 148586 429338 148822 429574
rect 148266 389658 148502 389894
rect 148586 389658 148822 389894
rect 148266 389338 148502 389574
rect 148586 389338 148822 389574
rect 148266 349658 148502 349894
rect 148586 349658 148822 349894
rect 148266 349338 148502 349574
rect 148586 349338 148822 349574
rect 148266 309658 148502 309894
rect 148586 309658 148822 309894
rect 148266 309338 148502 309574
rect 148586 309338 148822 309574
rect 148266 269658 148502 269894
rect 148586 269658 148822 269894
rect 148266 269338 148502 269574
rect 148586 269338 148822 269574
rect 148266 229658 148502 229894
rect 148586 229658 148822 229894
rect 148266 229338 148502 229574
rect 148586 229338 148822 229574
rect 148266 189658 148502 189894
rect 148586 189658 148822 189894
rect 148266 189338 148502 189574
rect 148586 189338 148822 189574
rect 148266 149658 148502 149894
rect 148586 149658 148822 149894
rect 148266 149338 148502 149574
rect 148586 149338 148822 149574
rect 148266 109658 148502 109894
rect 148586 109658 148822 109894
rect 148266 109338 148502 109574
rect 148586 109338 148822 109574
rect 148266 69658 148502 69894
rect 148586 69658 148822 69894
rect 148266 69338 148502 69574
rect 148586 69338 148822 69574
rect 148266 29658 148502 29894
rect 148586 29658 148822 29894
rect 148266 29338 148502 29574
rect 148586 29338 148822 29574
rect 148266 -5382 148502 -5146
rect 148586 -5382 148822 -5146
rect 148266 -5702 148502 -5466
rect 148586 -5702 148822 -5466
rect 171986 710362 172222 710598
rect 172306 710362 172542 710598
rect 171986 710042 172222 710278
rect 172306 710042 172542 710278
rect 168266 708442 168502 708678
rect 168586 708442 168822 708678
rect 168266 708122 168502 708358
rect 168586 708122 168822 708358
rect 164546 706522 164782 706758
rect 164866 706522 165102 706758
rect 164546 706202 164782 706438
rect 164866 706202 165102 706438
rect 151986 673378 152222 673614
rect 152306 673378 152542 673614
rect 151986 673058 152222 673294
rect 152306 673058 152542 673294
rect 151986 633378 152222 633614
rect 152306 633378 152542 633614
rect 151986 633058 152222 633294
rect 152306 633058 152542 633294
rect 151986 593378 152222 593614
rect 152306 593378 152542 593614
rect 151986 593058 152222 593294
rect 152306 593058 152542 593294
rect 151986 553378 152222 553614
rect 152306 553378 152542 553614
rect 151986 553058 152222 553294
rect 152306 553058 152542 553294
rect 151986 513378 152222 513614
rect 152306 513378 152542 513614
rect 151986 513058 152222 513294
rect 152306 513058 152542 513294
rect 151986 473378 152222 473614
rect 152306 473378 152542 473614
rect 151986 473058 152222 473294
rect 152306 473058 152542 473294
rect 151986 433378 152222 433614
rect 152306 433378 152542 433614
rect 151986 433058 152222 433294
rect 152306 433058 152542 433294
rect 151986 393378 152222 393614
rect 152306 393378 152542 393614
rect 151986 393058 152222 393294
rect 152306 393058 152542 393294
rect 151986 353378 152222 353614
rect 152306 353378 152542 353614
rect 151986 353058 152222 353294
rect 152306 353058 152542 353294
rect 160826 704602 161062 704838
rect 161146 704602 161382 704838
rect 160826 704282 161062 704518
rect 161146 704282 161382 704518
rect 160826 682218 161062 682454
rect 161146 682218 161382 682454
rect 160826 681898 161062 682134
rect 161146 681898 161382 682134
rect 160826 642218 161062 642454
rect 161146 642218 161382 642454
rect 160826 641898 161062 642134
rect 161146 641898 161382 642134
rect 160826 602218 161062 602454
rect 161146 602218 161382 602454
rect 160826 601898 161062 602134
rect 161146 601898 161382 602134
rect 160826 562218 161062 562454
rect 161146 562218 161382 562454
rect 160826 561898 161062 562134
rect 161146 561898 161382 562134
rect 160826 522218 161062 522454
rect 161146 522218 161382 522454
rect 160826 521898 161062 522134
rect 161146 521898 161382 522134
rect 160826 482218 161062 482454
rect 161146 482218 161382 482454
rect 160826 481898 161062 482134
rect 161146 481898 161382 482134
rect 160826 442218 161062 442454
rect 161146 442218 161382 442454
rect 160826 441898 161062 442134
rect 161146 441898 161382 442134
rect 160826 402218 161062 402454
rect 161146 402218 161382 402454
rect 160826 401898 161062 402134
rect 161146 401898 161382 402134
rect 160826 362218 161062 362454
rect 161146 362218 161382 362454
rect 160826 361898 161062 362134
rect 161146 361898 161382 362134
rect 160826 322218 161062 322454
rect 161146 322218 161382 322454
rect 160826 321898 161062 322134
rect 161146 321898 161382 322134
rect 151986 313378 152222 313614
rect 152306 313378 152542 313614
rect 151986 313058 152222 313294
rect 152306 313058 152542 313294
rect 151986 273378 152222 273614
rect 152306 273378 152542 273614
rect 151986 273058 152222 273294
rect 152306 273058 152542 273294
rect 151986 233378 152222 233614
rect 152306 233378 152542 233614
rect 151986 233058 152222 233294
rect 152306 233058 152542 233294
rect 151986 193378 152222 193614
rect 152306 193378 152542 193614
rect 151986 193058 152222 193294
rect 152306 193058 152542 193294
rect 151986 153378 152222 153614
rect 152306 153378 152542 153614
rect 151986 153058 152222 153294
rect 152306 153058 152542 153294
rect 151986 113378 152222 113614
rect 152306 113378 152542 113614
rect 151986 113058 152222 113294
rect 152306 113058 152542 113294
rect 151986 73378 152222 73614
rect 152306 73378 152542 73614
rect 151986 73058 152222 73294
rect 152306 73058 152542 73294
rect 151986 33378 152222 33614
rect 152306 33378 152542 33614
rect 151986 33058 152222 33294
rect 152306 33058 152542 33294
rect 131986 -6342 132222 -6106
rect 132306 -6342 132542 -6106
rect 131986 -6662 132222 -6426
rect 132306 -6662 132542 -6426
rect 160826 282218 161382 282454
rect 160826 281898 161382 282134
rect 160826 242218 161382 242454
rect 160826 241898 161382 242134
rect 160826 202218 161382 202454
rect 160826 201898 161382 202134
rect 160826 162218 161382 162454
rect 160826 161898 161382 162134
rect 160826 122218 161062 122454
rect 161146 122218 161382 122454
rect 160826 121898 161062 122134
rect 161146 121898 161382 122134
rect 160826 82218 161062 82454
rect 161146 82218 161382 82454
rect 160826 81898 161062 82134
rect 161146 81898 161382 82134
rect 160826 42218 161062 42454
rect 161146 42218 161382 42454
rect 160826 41898 161062 42134
rect 161146 41898 161382 42134
rect 160826 2218 161062 2454
rect 161146 2218 161382 2454
rect 160826 1898 161062 2134
rect 161146 1898 161382 2134
rect 160826 -582 161062 -346
rect 161146 -582 161382 -346
rect 160826 -902 161062 -666
rect 161146 -902 161382 -666
rect 164546 685938 164782 686174
rect 164866 685938 165102 686174
rect 164546 685618 164782 685854
rect 164866 685618 165102 685854
rect 164546 645938 164782 646174
rect 164866 645938 165102 646174
rect 164546 645618 164782 645854
rect 164866 645618 165102 645854
rect 164546 605938 164782 606174
rect 164866 605938 165102 606174
rect 164546 605618 164782 605854
rect 164866 605618 165102 605854
rect 164546 565938 164782 566174
rect 164866 565938 165102 566174
rect 164546 565618 164782 565854
rect 164866 565618 165102 565854
rect 164546 525938 164782 526174
rect 164866 525938 165102 526174
rect 164546 525618 164782 525854
rect 164866 525618 165102 525854
rect 164546 485938 164782 486174
rect 164866 485938 165102 486174
rect 164546 485618 164782 485854
rect 164866 485618 165102 485854
rect 164546 445938 164782 446174
rect 164866 445938 165102 446174
rect 164546 445618 164782 445854
rect 164866 445618 165102 445854
rect 164546 405938 164782 406174
rect 164866 405938 165102 406174
rect 164546 405618 164782 405854
rect 164866 405618 165102 405854
rect 164546 365938 164782 366174
rect 164866 365938 165102 366174
rect 164546 365618 164782 365854
rect 164866 365618 165102 365854
rect 164546 325938 164782 326174
rect 164866 325938 165102 326174
rect 164546 325618 164782 325854
rect 164866 325618 165102 325854
rect 164546 285938 164782 286174
rect 164866 285938 165102 286174
rect 164546 285618 164782 285854
rect 164866 285618 165102 285854
rect 164546 245938 164782 246174
rect 164866 245938 165102 246174
rect 164546 245618 164782 245854
rect 164866 245618 165102 245854
rect 164546 205938 164782 206174
rect 164866 205938 165102 206174
rect 164546 205618 164782 205854
rect 164866 205618 165102 205854
rect 164546 165938 164782 166174
rect 164866 165938 165102 166174
rect 164546 165618 164782 165854
rect 164866 165618 165102 165854
rect 164546 125938 164782 126174
rect 164866 125938 165102 126174
rect 164546 125618 164782 125854
rect 164866 125618 165102 125854
rect 164546 85938 164782 86174
rect 164866 85938 165102 86174
rect 164546 85618 164782 85854
rect 164866 85618 165102 85854
rect 164546 45938 164782 46174
rect 164866 45938 165102 46174
rect 164546 45618 164782 45854
rect 164866 45618 165102 45854
rect 164546 5938 164782 6174
rect 164866 5938 165102 6174
rect 164546 5618 164782 5854
rect 164866 5618 165102 5854
rect 164546 -2502 164782 -2266
rect 164866 -2502 165102 -2266
rect 164546 -2822 164782 -2586
rect 164866 -2822 165102 -2586
rect 168266 689658 168502 689894
rect 168586 689658 168822 689894
rect 168266 689338 168502 689574
rect 168586 689338 168822 689574
rect 168266 649658 168502 649894
rect 168586 649658 168822 649894
rect 168266 649338 168502 649574
rect 168586 649338 168822 649574
rect 168266 609658 168502 609894
rect 168586 609658 168822 609894
rect 168266 609338 168502 609574
rect 168586 609338 168822 609574
rect 168266 569658 168502 569894
rect 168586 569658 168822 569894
rect 168266 569338 168502 569574
rect 168586 569338 168822 569574
rect 168266 529658 168502 529894
rect 168586 529658 168822 529894
rect 168266 529338 168502 529574
rect 168586 529338 168822 529574
rect 168266 489658 168502 489894
rect 168586 489658 168822 489894
rect 168266 489338 168502 489574
rect 168586 489338 168822 489574
rect 168266 449658 168502 449894
rect 168586 449658 168822 449894
rect 168266 449338 168502 449574
rect 168586 449338 168822 449574
rect 168266 409658 168502 409894
rect 168586 409658 168822 409894
rect 168266 409338 168502 409574
rect 168586 409338 168822 409574
rect 168266 369658 168502 369894
rect 168586 369658 168822 369894
rect 168266 369338 168502 369574
rect 168586 369338 168822 369574
rect 168266 329658 168502 329894
rect 168586 329658 168822 329894
rect 168266 329338 168502 329574
rect 168586 329338 168822 329574
rect 191986 711322 192222 711558
rect 192306 711322 192542 711558
rect 191986 711002 192222 711238
rect 192306 711002 192542 711238
rect 188266 709402 188502 709638
rect 188586 709402 188822 709638
rect 188266 709082 188502 709318
rect 188586 709082 188822 709318
rect 184546 707482 184782 707718
rect 184866 707482 185102 707718
rect 184546 707162 184782 707398
rect 184866 707162 185102 707398
rect 171986 693378 172222 693614
rect 172306 693378 172542 693614
rect 171986 693058 172222 693294
rect 172306 693058 172542 693294
rect 171986 653378 172222 653614
rect 172306 653378 172542 653614
rect 171986 653058 172222 653294
rect 172306 653058 172542 653294
rect 171986 613378 172222 613614
rect 172306 613378 172542 613614
rect 171986 613058 172222 613294
rect 172306 613058 172542 613294
rect 171986 573378 172222 573614
rect 172306 573378 172542 573614
rect 171986 573058 172222 573294
rect 172306 573058 172542 573294
rect 171986 533378 172222 533614
rect 172306 533378 172542 533614
rect 171986 533058 172222 533294
rect 172306 533058 172542 533294
rect 171986 493378 172222 493614
rect 172306 493378 172542 493614
rect 171986 493058 172222 493294
rect 172306 493058 172542 493294
rect 171986 453378 172222 453614
rect 172306 453378 172542 453614
rect 171986 453058 172222 453294
rect 172306 453058 172542 453294
rect 171986 413378 172222 413614
rect 172306 413378 172542 413614
rect 171986 413058 172222 413294
rect 172306 413058 172542 413294
rect 171986 373378 172222 373614
rect 172306 373378 172542 373614
rect 171986 373058 172222 373294
rect 172306 373058 172542 373294
rect 171986 333378 172222 333614
rect 172306 333378 172542 333614
rect 171986 333058 172222 333294
rect 172306 333058 172542 333294
rect 168266 289658 168502 289894
rect 168586 289658 168822 289894
rect 168266 289338 168502 289574
rect 168586 289338 168822 289574
rect 168266 249658 168502 249894
rect 168586 249658 168822 249894
rect 168266 249338 168502 249574
rect 168586 249338 168822 249574
rect 168266 209658 168502 209894
rect 168586 209658 168822 209894
rect 168266 209338 168502 209574
rect 168586 209338 168822 209574
rect 168266 169658 168502 169894
rect 168586 169658 168822 169894
rect 168266 169338 168502 169574
rect 168586 169338 168822 169574
rect 168266 129658 168502 129894
rect 168586 129658 168822 129894
rect 168266 129338 168502 129574
rect 168586 129338 168822 129574
rect 168266 89658 168502 89894
rect 168586 89658 168822 89894
rect 168266 89338 168502 89574
rect 168586 89338 168822 89574
rect 168266 49658 168502 49894
rect 168586 49658 168822 49894
rect 168266 49338 168502 49574
rect 168586 49338 168822 49574
rect 168266 9658 168502 9894
rect 168586 9658 168822 9894
rect 168266 9338 168502 9574
rect 168586 9338 168822 9574
rect 180826 705562 181062 705798
rect 181146 705562 181382 705798
rect 180826 705242 181062 705478
rect 181146 705242 181382 705478
rect 180826 662218 181062 662454
rect 181146 662218 181382 662454
rect 180826 661898 181062 662134
rect 181146 661898 181382 662134
rect 180826 622218 181062 622454
rect 181146 622218 181382 622454
rect 180826 621898 181062 622134
rect 181146 621898 181382 622134
rect 180826 582218 181062 582454
rect 181146 582218 181382 582454
rect 180826 581898 181062 582134
rect 181146 581898 181382 582134
rect 180826 542218 181062 542454
rect 181146 542218 181382 542454
rect 180826 541898 181062 542134
rect 181146 541898 181382 542134
rect 180826 502218 181062 502454
rect 181146 502218 181382 502454
rect 180826 501898 181062 502134
rect 181146 501898 181382 502134
rect 180826 462218 181062 462454
rect 181146 462218 181382 462454
rect 180826 461898 181062 462134
rect 181146 461898 181382 462134
rect 180826 422218 181062 422454
rect 181146 422218 181382 422454
rect 180826 421898 181062 422134
rect 181146 421898 181382 422134
rect 180826 382218 181062 382454
rect 181146 382218 181382 382454
rect 180826 381898 181062 382134
rect 181146 381898 181382 382134
rect 180826 342218 181062 342454
rect 181146 342218 181382 342454
rect 180826 341898 181062 342134
rect 181146 341898 181382 342134
rect 171986 293378 172222 293614
rect 172306 293378 172542 293614
rect 171986 293058 172222 293294
rect 172306 293058 172542 293294
rect 171986 253378 172222 253614
rect 172306 253378 172542 253614
rect 171986 253058 172222 253294
rect 172306 253058 172542 253294
rect 171986 213378 172222 213614
rect 172306 213378 172542 213614
rect 171986 213058 172222 213294
rect 172306 213058 172542 213294
rect 171986 173378 172222 173614
rect 172306 173378 172542 173614
rect 171986 173058 172222 173294
rect 172306 173058 172542 173294
rect 171986 133378 172222 133614
rect 172306 133378 172542 133614
rect 171986 133058 172222 133294
rect 172306 133058 172542 133294
rect 171986 93378 172222 93614
rect 172306 93378 172542 93614
rect 171986 93058 172222 93294
rect 172306 93058 172542 93294
rect 171986 53378 172222 53614
rect 172306 53378 172542 53614
rect 171986 53058 172222 53294
rect 172306 53058 172542 53294
rect 171986 13378 172222 13614
rect 172306 13378 172542 13614
rect 171986 13058 172222 13294
rect 172306 13058 172542 13294
rect 168266 -4422 168502 -4186
rect 168586 -4422 168822 -4186
rect 168266 -4742 168502 -4506
rect 168586 -4742 168822 -4506
rect 151986 -7302 152222 -7066
rect 152306 -7302 152542 -7066
rect 151986 -7622 152222 -7386
rect 152306 -7622 152542 -7386
rect 180826 302218 181382 302454
rect 180826 301898 181382 302134
rect 180826 262218 181382 262454
rect 180826 261898 181382 262134
rect 180826 222218 181382 222454
rect 180826 221898 181382 222134
rect 180826 182218 181382 182454
rect 180826 181898 181382 182134
rect 180826 142218 181382 142454
rect 180826 141898 181382 142134
rect 180826 102218 181062 102454
rect 181146 102218 181382 102454
rect 180826 101898 181062 102134
rect 181146 101898 181382 102134
rect 180826 62218 181062 62454
rect 181146 62218 181382 62454
rect 180826 61898 181062 62134
rect 181146 61898 181382 62134
rect 180826 22218 181062 22454
rect 181146 22218 181382 22454
rect 180826 21898 181062 22134
rect 181146 21898 181382 22134
rect 180826 -1542 181062 -1306
rect 181146 -1542 181382 -1306
rect 180826 -1862 181062 -1626
rect 181146 -1862 181382 -1626
rect 184546 665938 184782 666174
rect 184866 665938 185102 666174
rect 184546 665618 184782 665854
rect 184866 665618 185102 665854
rect 184546 625938 184782 626174
rect 184866 625938 185102 626174
rect 184546 625618 184782 625854
rect 184866 625618 185102 625854
rect 184546 585938 184782 586174
rect 184866 585938 185102 586174
rect 184546 585618 184782 585854
rect 184866 585618 185102 585854
rect 184546 545938 184782 546174
rect 184866 545938 185102 546174
rect 184546 545618 184782 545854
rect 184866 545618 185102 545854
rect 184546 505938 184782 506174
rect 184866 505938 185102 506174
rect 184546 505618 184782 505854
rect 184866 505618 185102 505854
rect 184546 465938 184782 466174
rect 184866 465938 185102 466174
rect 184546 465618 184782 465854
rect 184866 465618 185102 465854
rect 184546 425938 184782 426174
rect 184866 425938 185102 426174
rect 184546 425618 184782 425854
rect 184866 425618 185102 425854
rect 184546 385938 184782 386174
rect 184866 385938 185102 386174
rect 184546 385618 184782 385854
rect 184866 385618 185102 385854
rect 184546 345938 184782 346174
rect 184866 345938 185102 346174
rect 184546 345618 184782 345854
rect 184866 345618 185102 345854
rect 184546 305938 184782 306174
rect 184866 305938 185102 306174
rect 184546 305618 184782 305854
rect 184866 305618 185102 305854
rect 184546 265938 184782 266174
rect 184866 265938 185102 266174
rect 184546 265618 184782 265854
rect 184866 265618 185102 265854
rect 184546 225938 184782 226174
rect 184866 225938 185102 226174
rect 184546 225618 184782 225854
rect 184866 225618 185102 225854
rect 184546 185938 184782 186174
rect 184866 185938 185102 186174
rect 184546 185618 184782 185854
rect 184866 185618 185102 185854
rect 184546 145938 184782 146174
rect 184866 145938 185102 146174
rect 184546 145618 184782 145854
rect 184866 145618 185102 145854
rect 184546 105938 184782 106174
rect 184866 105938 185102 106174
rect 184546 105618 184782 105854
rect 184866 105618 185102 105854
rect 184546 65938 184782 66174
rect 184866 65938 185102 66174
rect 184546 65618 184782 65854
rect 184866 65618 185102 65854
rect 184546 25938 184782 26174
rect 184866 25938 185102 26174
rect 184546 25618 184782 25854
rect 184866 25618 185102 25854
rect 184546 -3462 184782 -3226
rect 184866 -3462 185102 -3226
rect 184546 -3782 184782 -3546
rect 184866 -3782 185102 -3546
rect 188266 669658 188502 669894
rect 188586 669658 188822 669894
rect 188266 669338 188502 669574
rect 188586 669338 188822 669574
rect 188266 629658 188502 629894
rect 188586 629658 188822 629894
rect 188266 629338 188502 629574
rect 188586 629338 188822 629574
rect 188266 589658 188502 589894
rect 188586 589658 188822 589894
rect 188266 589338 188502 589574
rect 188586 589338 188822 589574
rect 188266 549658 188502 549894
rect 188586 549658 188822 549894
rect 188266 549338 188502 549574
rect 188586 549338 188822 549574
rect 188266 509658 188502 509894
rect 188586 509658 188822 509894
rect 188266 509338 188502 509574
rect 188586 509338 188822 509574
rect 188266 469658 188502 469894
rect 188586 469658 188822 469894
rect 188266 469338 188502 469574
rect 188586 469338 188822 469574
rect 188266 429658 188502 429894
rect 188586 429658 188822 429894
rect 188266 429338 188502 429574
rect 188586 429338 188822 429574
rect 188266 389658 188502 389894
rect 188586 389658 188822 389894
rect 188266 389338 188502 389574
rect 188586 389338 188822 389574
rect 188266 349658 188502 349894
rect 188586 349658 188822 349894
rect 188266 349338 188502 349574
rect 188586 349338 188822 349574
rect 188266 309658 188502 309894
rect 188586 309658 188822 309894
rect 188266 309338 188502 309574
rect 188586 309338 188822 309574
rect 188266 269658 188502 269894
rect 188586 269658 188822 269894
rect 188266 269338 188502 269574
rect 188586 269338 188822 269574
rect 188266 229658 188502 229894
rect 188586 229658 188822 229894
rect 188266 229338 188502 229574
rect 188586 229338 188822 229574
rect 188266 189658 188502 189894
rect 188586 189658 188822 189894
rect 188266 189338 188502 189574
rect 188586 189338 188822 189574
rect 188266 149658 188502 149894
rect 188586 149658 188822 149894
rect 188266 149338 188502 149574
rect 188586 149338 188822 149574
rect 188266 109658 188502 109894
rect 188586 109658 188822 109894
rect 188266 109338 188502 109574
rect 188586 109338 188822 109574
rect 188266 69658 188502 69894
rect 188586 69658 188822 69894
rect 188266 69338 188502 69574
rect 188586 69338 188822 69574
rect 188266 29658 188502 29894
rect 188586 29658 188822 29894
rect 188266 29338 188502 29574
rect 188586 29338 188822 29574
rect 188266 -5382 188502 -5146
rect 188586 -5382 188822 -5146
rect 188266 -5702 188502 -5466
rect 188586 -5702 188822 -5466
rect 211986 710362 212222 710598
rect 212306 710362 212542 710598
rect 211986 710042 212222 710278
rect 212306 710042 212542 710278
rect 208266 708442 208502 708678
rect 208586 708442 208822 708678
rect 208266 708122 208502 708358
rect 208586 708122 208822 708358
rect 204546 706522 204782 706758
rect 204866 706522 205102 706758
rect 204546 706202 204782 706438
rect 204866 706202 205102 706438
rect 191986 673378 192222 673614
rect 192306 673378 192542 673614
rect 191986 673058 192222 673294
rect 192306 673058 192542 673294
rect 191986 633378 192222 633614
rect 192306 633378 192542 633614
rect 191986 633058 192222 633294
rect 192306 633058 192542 633294
rect 191986 593378 192222 593614
rect 192306 593378 192542 593614
rect 191986 593058 192222 593294
rect 192306 593058 192542 593294
rect 191986 553378 192222 553614
rect 192306 553378 192542 553614
rect 191986 553058 192222 553294
rect 192306 553058 192542 553294
rect 191986 513378 192222 513614
rect 192306 513378 192542 513614
rect 191986 513058 192222 513294
rect 192306 513058 192542 513294
rect 191986 473378 192222 473614
rect 192306 473378 192542 473614
rect 191986 473058 192222 473294
rect 192306 473058 192542 473294
rect 191986 433378 192222 433614
rect 192306 433378 192542 433614
rect 191986 433058 192222 433294
rect 192306 433058 192542 433294
rect 191986 393378 192222 393614
rect 192306 393378 192542 393614
rect 191986 393058 192222 393294
rect 192306 393058 192542 393294
rect 191986 353378 192222 353614
rect 192306 353378 192542 353614
rect 191986 353058 192222 353294
rect 192306 353058 192542 353294
rect 200826 704602 201062 704838
rect 201146 704602 201382 704838
rect 200826 704282 201062 704518
rect 201146 704282 201382 704518
rect 200826 682218 201062 682454
rect 201146 682218 201382 682454
rect 200826 681898 201062 682134
rect 201146 681898 201382 682134
rect 200826 642218 201062 642454
rect 201146 642218 201382 642454
rect 200826 641898 201062 642134
rect 201146 641898 201382 642134
rect 200826 602218 201062 602454
rect 201146 602218 201382 602454
rect 200826 601898 201062 602134
rect 201146 601898 201382 602134
rect 200826 562218 201062 562454
rect 201146 562218 201382 562454
rect 200826 561898 201062 562134
rect 201146 561898 201382 562134
rect 200826 522218 201062 522454
rect 201146 522218 201382 522454
rect 200826 521898 201062 522134
rect 201146 521898 201382 522134
rect 200826 482218 201062 482454
rect 201146 482218 201382 482454
rect 200826 481898 201062 482134
rect 201146 481898 201382 482134
rect 200826 442218 201062 442454
rect 201146 442218 201382 442454
rect 200826 441898 201062 442134
rect 201146 441898 201382 442134
rect 200826 402218 201062 402454
rect 201146 402218 201382 402454
rect 200826 401898 201062 402134
rect 201146 401898 201382 402134
rect 200826 362218 201062 362454
rect 201146 362218 201382 362454
rect 200826 361898 201062 362134
rect 201146 361898 201382 362134
rect 200826 322218 201062 322454
rect 201146 322218 201382 322454
rect 200826 321898 201062 322134
rect 201146 321898 201382 322134
rect 191986 313378 192222 313614
rect 192306 313378 192542 313614
rect 191986 313058 192222 313294
rect 192306 313058 192542 313294
rect 191986 273378 192222 273614
rect 192306 273378 192542 273614
rect 191986 273058 192222 273294
rect 192306 273058 192542 273294
rect 191986 233378 192222 233614
rect 192306 233378 192542 233614
rect 191986 233058 192222 233294
rect 192306 233058 192542 233294
rect 191986 193378 192222 193614
rect 192306 193378 192542 193614
rect 191986 193058 192222 193294
rect 192306 193058 192542 193294
rect 191986 153378 192222 153614
rect 192306 153378 192542 153614
rect 191986 153058 192222 153294
rect 192306 153058 192542 153294
rect 191986 113378 192222 113614
rect 192306 113378 192542 113614
rect 191986 113058 192222 113294
rect 192306 113058 192542 113294
rect 191986 73378 192222 73614
rect 192306 73378 192542 73614
rect 191986 73058 192222 73294
rect 192306 73058 192542 73294
rect 191986 33378 192222 33614
rect 192306 33378 192542 33614
rect 191986 33058 192222 33294
rect 192306 33058 192542 33294
rect 171986 -6342 172222 -6106
rect 172306 -6342 172542 -6106
rect 171986 -6662 172222 -6426
rect 172306 -6662 172542 -6426
rect 200826 282218 201382 282454
rect 200826 281898 201382 282134
rect 200826 242218 201382 242454
rect 200826 241898 201382 242134
rect 200826 202218 201382 202454
rect 200826 201898 201382 202134
rect 200826 162218 201382 162454
rect 200826 161898 201382 162134
rect 200826 122218 201062 122454
rect 201146 122218 201382 122454
rect 200826 121898 201062 122134
rect 201146 121898 201382 122134
rect 200826 82218 201062 82454
rect 201146 82218 201382 82454
rect 200826 81898 201062 82134
rect 201146 81898 201382 82134
rect 200826 42218 201062 42454
rect 201146 42218 201382 42454
rect 200826 41898 201062 42134
rect 201146 41898 201382 42134
rect 200826 2218 201062 2454
rect 201146 2218 201382 2454
rect 200826 1898 201062 2134
rect 201146 1898 201382 2134
rect 200826 -582 201062 -346
rect 201146 -582 201382 -346
rect 200826 -902 201062 -666
rect 201146 -902 201382 -666
rect 204546 685938 204782 686174
rect 204866 685938 205102 686174
rect 204546 685618 204782 685854
rect 204866 685618 205102 685854
rect 204546 645938 204782 646174
rect 204866 645938 205102 646174
rect 204546 645618 204782 645854
rect 204866 645618 205102 645854
rect 204546 605938 204782 606174
rect 204866 605938 205102 606174
rect 204546 605618 204782 605854
rect 204866 605618 205102 605854
rect 204546 565938 204782 566174
rect 204866 565938 205102 566174
rect 204546 565618 204782 565854
rect 204866 565618 205102 565854
rect 204546 525938 204782 526174
rect 204866 525938 205102 526174
rect 204546 525618 204782 525854
rect 204866 525618 205102 525854
rect 204546 485938 204782 486174
rect 204866 485938 205102 486174
rect 204546 485618 204782 485854
rect 204866 485618 205102 485854
rect 204546 445938 204782 446174
rect 204866 445938 205102 446174
rect 204546 445618 204782 445854
rect 204866 445618 205102 445854
rect 204546 405938 204782 406174
rect 204866 405938 205102 406174
rect 204546 405618 204782 405854
rect 204866 405618 205102 405854
rect 204546 365938 204782 366174
rect 204866 365938 205102 366174
rect 204546 365618 204782 365854
rect 204866 365618 205102 365854
rect 204546 325938 204782 326174
rect 204866 325938 205102 326174
rect 204546 325618 204782 325854
rect 204866 325618 205102 325854
rect 204546 285938 204782 286174
rect 204866 285938 205102 286174
rect 204546 285618 204782 285854
rect 204866 285618 205102 285854
rect 204546 245938 204782 246174
rect 204866 245938 205102 246174
rect 204546 245618 204782 245854
rect 204866 245618 205102 245854
rect 204546 205938 204782 206174
rect 204866 205938 205102 206174
rect 204546 205618 204782 205854
rect 204866 205618 205102 205854
rect 204546 165938 204782 166174
rect 204866 165938 205102 166174
rect 204546 165618 204782 165854
rect 204866 165618 205102 165854
rect 204546 125938 204782 126174
rect 204866 125938 205102 126174
rect 204546 125618 204782 125854
rect 204866 125618 205102 125854
rect 204546 85938 204782 86174
rect 204866 85938 205102 86174
rect 204546 85618 204782 85854
rect 204866 85618 205102 85854
rect 204546 45938 204782 46174
rect 204866 45938 205102 46174
rect 204546 45618 204782 45854
rect 204866 45618 205102 45854
rect 204546 5938 204782 6174
rect 204866 5938 205102 6174
rect 204546 5618 204782 5854
rect 204866 5618 205102 5854
rect 204546 -2502 204782 -2266
rect 204866 -2502 205102 -2266
rect 204546 -2822 204782 -2586
rect 204866 -2822 205102 -2586
rect 208266 689658 208502 689894
rect 208586 689658 208822 689894
rect 208266 689338 208502 689574
rect 208586 689338 208822 689574
rect 208266 649658 208502 649894
rect 208586 649658 208822 649894
rect 208266 649338 208502 649574
rect 208586 649338 208822 649574
rect 208266 609658 208502 609894
rect 208586 609658 208822 609894
rect 208266 609338 208502 609574
rect 208586 609338 208822 609574
rect 208266 569658 208502 569894
rect 208586 569658 208822 569894
rect 208266 569338 208502 569574
rect 208586 569338 208822 569574
rect 208266 529658 208502 529894
rect 208586 529658 208822 529894
rect 208266 529338 208502 529574
rect 208586 529338 208822 529574
rect 208266 489658 208502 489894
rect 208586 489658 208822 489894
rect 208266 489338 208502 489574
rect 208586 489338 208822 489574
rect 208266 449658 208502 449894
rect 208586 449658 208822 449894
rect 208266 449338 208502 449574
rect 208586 449338 208822 449574
rect 208266 409658 208502 409894
rect 208586 409658 208822 409894
rect 208266 409338 208502 409574
rect 208586 409338 208822 409574
rect 208266 369658 208502 369894
rect 208586 369658 208822 369894
rect 208266 369338 208502 369574
rect 208586 369338 208822 369574
rect 208266 329658 208502 329894
rect 208586 329658 208822 329894
rect 208266 329338 208502 329574
rect 208586 329338 208822 329574
rect 208266 289658 208502 289894
rect 208586 289658 208822 289894
rect 208266 289338 208502 289574
rect 208586 289338 208822 289574
rect 208266 249658 208502 249894
rect 208586 249658 208822 249894
rect 208266 249338 208502 249574
rect 208586 249338 208822 249574
rect 208266 209658 208502 209894
rect 208586 209658 208822 209894
rect 208266 209338 208502 209574
rect 208586 209338 208822 209574
rect 208266 169658 208502 169894
rect 208586 169658 208822 169894
rect 208266 169338 208502 169574
rect 208586 169338 208822 169574
rect 208266 129658 208502 129894
rect 208586 129658 208822 129894
rect 208266 129338 208502 129574
rect 208586 129338 208822 129574
rect 208266 89658 208502 89894
rect 208586 89658 208822 89894
rect 208266 89338 208502 89574
rect 208586 89338 208822 89574
rect 208266 49658 208502 49894
rect 208586 49658 208822 49894
rect 208266 49338 208502 49574
rect 208586 49338 208822 49574
rect 208266 9658 208502 9894
rect 208586 9658 208822 9894
rect 208266 9338 208502 9574
rect 208586 9338 208822 9574
rect 208266 -4422 208502 -4186
rect 208586 -4422 208822 -4186
rect 208266 -4742 208502 -4506
rect 208586 -4742 208822 -4506
rect 231986 711322 232222 711558
rect 232306 711322 232542 711558
rect 231986 711002 232222 711238
rect 232306 711002 232542 711238
rect 228266 709402 228502 709638
rect 228586 709402 228822 709638
rect 228266 709082 228502 709318
rect 228586 709082 228822 709318
rect 224546 707482 224782 707718
rect 224866 707482 225102 707718
rect 224546 707162 224782 707398
rect 224866 707162 225102 707398
rect 211986 693378 212222 693614
rect 212306 693378 212542 693614
rect 211986 693058 212222 693294
rect 212306 693058 212542 693294
rect 211986 653378 212222 653614
rect 212306 653378 212542 653614
rect 211986 653058 212222 653294
rect 212306 653058 212542 653294
rect 211986 613378 212222 613614
rect 212306 613378 212542 613614
rect 211986 613058 212222 613294
rect 212306 613058 212542 613294
rect 211986 573378 212222 573614
rect 212306 573378 212542 573614
rect 211986 573058 212222 573294
rect 212306 573058 212542 573294
rect 211986 533378 212222 533614
rect 212306 533378 212542 533614
rect 211986 533058 212222 533294
rect 212306 533058 212542 533294
rect 211986 493378 212222 493614
rect 212306 493378 212542 493614
rect 211986 493058 212222 493294
rect 212306 493058 212542 493294
rect 211986 453378 212222 453614
rect 212306 453378 212542 453614
rect 211986 453058 212222 453294
rect 212306 453058 212542 453294
rect 211986 413378 212222 413614
rect 212306 413378 212542 413614
rect 211986 413058 212222 413294
rect 212306 413058 212542 413294
rect 211986 373378 212222 373614
rect 212306 373378 212542 373614
rect 211986 373058 212222 373294
rect 212306 373058 212542 373294
rect 211986 333378 212222 333614
rect 212306 333378 212542 333614
rect 211986 333058 212222 333294
rect 212306 333058 212542 333294
rect 211986 293378 212222 293614
rect 212306 293378 212542 293614
rect 211986 293058 212222 293294
rect 212306 293058 212542 293294
rect 211986 253378 212222 253614
rect 212306 253378 212542 253614
rect 211986 253058 212222 253294
rect 212306 253058 212542 253294
rect 211986 213378 212222 213614
rect 212306 213378 212542 213614
rect 211986 213058 212222 213294
rect 212306 213058 212542 213294
rect 211986 173378 212222 173614
rect 212306 173378 212542 173614
rect 211986 173058 212222 173294
rect 212306 173058 212542 173294
rect 211986 133378 212222 133614
rect 212306 133378 212542 133614
rect 211986 133058 212222 133294
rect 212306 133058 212542 133294
rect 211986 93378 212222 93614
rect 212306 93378 212542 93614
rect 211986 93058 212222 93294
rect 212306 93058 212542 93294
rect 211986 53378 212222 53614
rect 212306 53378 212542 53614
rect 211986 53058 212222 53294
rect 212306 53058 212542 53294
rect 211986 13378 212222 13614
rect 212306 13378 212542 13614
rect 211986 13058 212222 13294
rect 212306 13058 212542 13294
rect 191986 -7302 192222 -7066
rect 192306 -7302 192542 -7066
rect 191986 -7622 192222 -7386
rect 192306 -7622 192542 -7386
rect 220826 705562 221062 705798
rect 221146 705562 221382 705798
rect 220826 705242 221062 705478
rect 221146 705242 221382 705478
rect 220826 662218 221062 662454
rect 221146 662218 221382 662454
rect 220826 661898 221062 662134
rect 221146 661898 221382 662134
rect 220826 622218 221062 622454
rect 221146 622218 221382 622454
rect 220826 621898 221062 622134
rect 221146 621898 221382 622134
rect 220826 582218 221062 582454
rect 221146 582218 221382 582454
rect 220826 581898 221062 582134
rect 221146 581898 221382 582134
rect 220826 542218 221062 542454
rect 221146 542218 221382 542454
rect 220826 541898 221062 542134
rect 221146 541898 221382 542134
rect 220826 502218 221062 502454
rect 221146 502218 221382 502454
rect 220826 501898 221062 502134
rect 221146 501898 221382 502134
rect 220826 462218 221062 462454
rect 221146 462218 221382 462454
rect 220826 461898 221062 462134
rect 221146 461898 221382 462134
rect 220826 422218 221062 422454
rect 221146 422218 221382 422454
rect 220826 421898 221062 422134
rect 221146 421898 221382 422134
rect 220826 382218 221062 382454
rect 221146 382218 221382 382454
rect 220826 381898 221062 382134
rect 221146 381898 221382 382134
rect 220826 342218 221062 342454
rect 221146 342218 221382 342454
rect 220826 341898 221062 342134
rect 221146 341898 221382 342134
rect 220826 302218 221382 302454
rect 220826 301898 221382 302134
rect 220826 262218 221382 262454
rect 220826 261898 221382 262134
rect 220826 222218 221382 222454
rect 220826 221898 221382 222134
rect 220826 182218 221382 182454
rect 220826 181898 221382 182134
rect 220826 142218 221382 142454
rect 220826 141898 221382 142134
rect 220826 102218 221062 102454
rect 221146 102218 221382 102454
rect 220826 101898 221062 102134
rect 221146 101898 221382 102134
rect 220826 62218 221062 62454
rect 221146 62218 221382 62454
rect 220826 61898 221062 62134
rect 221146 61898 221382 62134
rect 220826 22218 221062 22454
rect 221146 22218 221382 22454
rect 220826 21898 221062 22134
rect 221146 21898 221382 22134
rect 220826 -1542 221062 -1306
rect 221146 -1542 221382 -1306
rect 220826 -1862 221062 -1626
rect 221146 -1862 221382 -1626
rect 224546 665938 224782 666174
rect 224866 665938 225102 666174
rect 224546 665618 224782 665854
rect 224866 665618 225102 665854
rect 224546 625938 224782 626174
rect 224866 625938 225102 626174
rect 224546 625618 224782 625854
rect 224866 625618 225102 625854
rect 224546 585938 224782 586174
rect 224866 585938 225102 586174
rect 224546 585618 224782 585854
rect 224866 585618 225102 585854
rect 224546 545938 224782 546174
rect 224866 545938 225102 546174
rect 224546 545618 224782 545854
rect 224866 545618 225102 545854
rect 224546 505938 224782 506174
rect 224866 505938 225102 506174
rect 224546 505618 224782 505854
rect 224866 505618 225102 505854
rect 224546 465938 224782 466174
rect 224866 465938 225102 466174
rect 224546 465618 224782 465854
rect 224866 465618 225102 465854
rect 224546 425938 224782 426174
rect 224866 425938 225102 426174
rect 224546 425618 224782 425854
rect 224866 425618 225102 425854
rect 224546 385938 224782 386174
rect 224866 385938 225102 386174
rect 224546 385618 224782 385854
rect 224866 385618 225102 385854
rect 224546 345938 224782 346174
rect 224866 345938 225102 346174
rect 224546 345618 224782 345854
rect 224866 345618 225102 345854
rect 224546 305938 224782 306174
rect 224866 305938 225102 306174
rect 224546 305618 224782 305854
rect 224866 305618 225102 305854
rect 224546 265938 224782 266174
rect 224866 265938 225102 266174
rect 224546 265618 224782 265854
rect 224866 265618 225102 265854
rect 224546 225938 224782 226174
rect 224866 225938 225102 226174
rect 224546 225618 224782 225854
rect 224866 225618 225102 225854
rect 224546 185938 224782 186174
rect 224866 185938 225102 186174
rect 224546 185618 224782 185854
rect 224866 185618 225102 185854
rect 224546 145938 224782 146174
rect 224866 145938 225102 146174
rect 224546 145618 224782 145854
rect 224866 145618 225102 145854
rect 224546 105938 224782 106174
rect 224866 105938 225102 106174
rect 224546 105618 224782 105854
rect 224866 105618 225102 105854
rect 224546 65938 224782 66174
rect 224866 65938 225102 66174
rect 224546 65618 224782 65854
rect 224866 65618 225102 65854
rect 224546 25938 224782 26174
rect 224866 25938 225102 26174
rect 224546 25618 224782 25854
rect 224866 25618 225102 25854
rect 224546 -3462 224782 -3226
rect 224866 -3462 225102 -3226
rect 224546 -3782 224782 -3546
rect 224866 -3782 225102 -3546
rect 228266 669658 228502 669894
rect 228586 669658 228822 669894
rect 228266 669338 228502 669574
rect 228586 669338 228822 669574
rect 228266 629658 228502 629894
rect 228586 629658 228822 629894
rect 228266 629338 228502 629574
rect 228586 629338 228822 629574
rect 228266 589658 228502 589894
rect 228586 589658 228822 589894
rect 228266 589338 228502 589574
rect 228586 589338 228822 589574
rect 228266 549658 228502 549894
rect 228586 549658 228822 549894
rect 228266 549338 228502 549574
rect 228586 549338 228822 549574
rect 228266 509658 228502 509894
rect 228586 509658 228822 509894
rect 228266 509338 228502 509574
rect 228586 509338 228822 509574
rect 228266 469658 228502 469894
rect 228586 469658 228822 469894
rect 228266 469338 228502 469574
rect 228586 469338 228822 469574
rect 228266 429658 228502 429894
rect 228586 429658 228822 429894
rect 228266 429338 228502 429574
rect 228586 429338 228822 429574
rect 228266 389658 228502 389894
rect 228586 389658 228822 389894
rect 228266 389338 228502 389574
rect 228586 389338 228822 389574
rect 228266 349658 228502 349894
rect 228586 349658 228822 349894
rect 228266 349338 228502 349574
rect 228586 349338 228822 349574
rect 228266 309658 228502 309894
rect 228586 309658 228822 309894
rect 228266 309338 228502 309574
rect 228586 309338 228822 309574
rect 228266 269658 228502 269894
rect 228586 269658 228822 269894
rect 228266 269338 228502 269574
rect 228586 269338 228822 269574
rect 228266 229658 228502 229894
rect 228586 229658 228822 229894
rect 228266 229338 228502 229574
rect 228586 229338 228822 229574
rect 228266 189658 228502 189894
rect 228586 189658 228822 189894
rect 228266 189338 228502 189574
rect 228586 189338 228822 189574
rect 228266 149658 228502 149894
rect 228586 149658 228822 149894
rect 228266 149338 228502 149574
rect 228586 149338 228822 149574
rect 228266 109658 228502 109894
rect 228586 109658 228822 109894
rect 228266 109338 228502 109574
rect 228586 109338 228822 109574
rect 228266 69658 228502 69894
rect 228586 69658 228822 69894
rect 228266 69338 228502 69574
rect 228586 69338 228822 69574
rect 228266 29658 228502 29894
rect 228586 29658 228822 29894
rect 228266 29338 228502 29574
rect 228586 29338 228822 29574
rect 228266 -5382 228502 -5146
rect 228586 -5382 228822 -5146
rect 228266 -5702 228502 -5466
rect 228586 -5702 228822 -5466
rect 251986 710362 252222 710598
rect 252306 710362 252542 710598
rect 251986 710042 252222 710278
rect 252306 710042 252542 710278
rect 248266 708442 248502 708678
rect 248586 708442 248822 708678
rect 248266 708122 248502 708358
rect 248586 708122 248822 708358
rect 244546 706522 244782 706758
rect 244866 706522 245102 706758
rect 244546 706202 244782 706438
rect 244866 706202 245102 706438
rect 231986 673378 232222 673614
rect 232306 673378 232542 673614
rect 231986 673058 232222 673294
rect 232306 673058 232542 673294
rect 231986 633378 232222 633614
rect 232306 633378 232542 633614
rect 231986 633058 232222 633294
rect 232306 633058 232542 633294
rect 231986 593378 232222 593614
rect 232306 593378 232542 593614
rect 231986 593058 232222 593294
rect 232306 593058 232542 593294
rect 231986 553378 232222 553614
rect 232306 553378 232542 553614
rect 231986 553058 232222 553294
rect 232306 553058 232542 553294
rect 231986 513378 232222 513614
rect 232306 513378 232542 513614
rect 231986 513058 232222 513294
rect 232306 513058 232542 513294
rect 231986 473378 232222 473614
rect 232306 473378 232542 473614
rect 231986 473058 232222 473294
rect 232306 473058 232542 473294
rect 231986 433378 232222 433614
rect 232306 433378 232542 433614
rect 231986 433058 232222 433294
rect 232306 433058 232542 433294
rect 231986 393378 232222 393614
rect 232306 393378 232542 393614
rect 231986 393058 232222 393294
rect 232306 393058 232542 393294
rect 231986 353378 232222 353614
rect 232306 353378 232542 353614
rect 231986 353058 232222 353294
rect 232306 353058 232542 353294
rect 240826 704602 241062 704838
rect 241146 704602 241382 704838
rect 240826 704282 241062 704518
rect 241146 704282 241382 704518
rect 240826 682218 241062 682454
rect 241146 682218 241382 682454
rect 240826 681898 241062 682134
rect 241146 681898 241382 682134
rect 240826 642218 241062 642454
rect 241146 642218 241382 642454
rect 240826 641898 241062 642134
rect 241146 641898 241382 642134
rect 240826 602218 241062 602454
rect 241146 602218 241382 602454
rect 240826 601898 241062 602134
rect 241146 601898 241382 602134
rect 240826 562218 241062 562454
rect 241146 562218 241382 562454
rect 240826 561898 241062 562134
rect 241146 561898 241382 562134
rect 240826 522218 241062 522454
rect 241146 522218 241382 522454
rect 240826 521898 241062 522134
rect 241146 521898 241382 522134
rect 240826 482218 241062 482454
rect 241146 482218 241382 482454
rect 240826 481898 241062 482134
rect 241146 481898 241382 482134
rect 240826 442218 241062 442454
rect 241146 442218 241382 442454
rect 240826 441898 241062 442134
rect 241146 441898 241382 442134
rect 240826 402218 241062 402454
rect 241146 402218 241382 402454
rect 240826 401898 241062 402134
rect 241146 401898 241382 402134
rect 240826 362218 241062 362454
rect 241146 362218 241382 362454
rect 240826 361898 241062 362134
rect 241146 361898 241382 362134
rect 240826 322218 241062 322454
rect 241146 322218 241382 322454
rect 240826 321898 241062 322134
rect 241146 321898 241382 322134
rect 231986 313378 232222 313614
rect 232306 313378 232542 313614
rect 231986 313058 232222 313294
rect 232306 313058 232542 313294
rect 231986 273378 232222 273614
rect 232306 273378 232542 273614
rect 231986 273058 232222 273294
rect 232306 273058 232542 273294
rect 231986 233378 232222 233614
rect 232306 233378 232542 233614
rect 231986 233058 232222 233294
rect 232306 233058 232542 233294
rect 231986 193378 232222 193614
rect 232306 193378 232542 193614
rect 231986 193058 232222 193294
rect 232306 193058 232542 193294
rect 231986 153378 232222 153614
rect 232306 153378 232542 153614
rect 231986 153058 232222 153294
rect 232306 153058 232542 153294
rect 231986 113378 232222 113614
rect 232306 113378 232542 113614
rect 231986 113058 232222 113294
rect 232306 113058 232542 113294
rect 231986 73378 232222 73614
rect 232306 73378 232542 73614
rect 231986 73058 232222 73294
rect 232306 73058 232542 73294
rect 231986 33378 232222 33614
rect 232306 33378 232542 33614
rect 231986 33058 232222 33294
rect 232306 33058 232542 33294
rect 211986 -6342 212222 -6106
rect 212306 -6342 212542 -6106
rect 211986 -6662 212222 -6426
rect 212306 -6662 212542 -6426
rect 240826 282218 241382 282454
rect 240826 281898 241382 282134
rect 240826 242218 241382 242454
rect 240826 241898 241382 242134
rect 240826 202218 241382 202454
rect 240826 201898 241382 202134
rect 240826 162218 241382 162454
rect 240826 161898 241382 162134
rect 240826 122218 241062 122454
rect 241146 122218 241382 122454
rect 240826 121898 241062 122134
rect 241146 121898 241382 122134
rect 240826 82218 241062 82454
rect 241146 82218 241382 82454
rect 240826 81898 241062 82134
rect 241146 81898 241382 82134
rect 240826 42218 241062 42454
rect 241146 42218 241382 42454
rect 240826 41898 241062 42134
rect 241146 41898 241382 42134
rect 240826 2218 241062 2454
rect 241146 2218 241382 2454
rect 240826 1898 241062 2134
rect 241146 1898 241382 2134
rect 240826 -582 241062 -346
rect 241146 -582 241382 -346
rect 240826 -902 241062 -666
rect 241146 -902 241382 -666
rect 244546 685938 244782 686174
rect 244866 685938 245102 686174
rect 244546 685618 244782 685854
rect 244866 685618 245102 685854
rect 244546 645938 244782 646174
rect 244866 645938 245102 646174
rect 244546 645618 244782 645854
rect 244866 645618 245102 645854
rect 244546 605938 244782 606174
rect 244866 605938 245102 606174
rect 244546 605618 244782 605854
rect 244866 605618 245102 605854
rect 244546 565938 244782 566174
rect 244866 565938 245102 566174
rect 244546 565618 244782 565854
rect 244866 565618 245102 565854
rect 244546 525938 244782 526174
rect 244866 525938 245102 526174
rect 244546 525618 244782 525854
rect 244866 525618 245102 525854
rect 244546 485938 244782 486174
rect 244866 485938 245102 486174
rect 244546 485618 244782 485854
rect 244866 485618 245102 485854
rect 244546 445938 244782 446174
rect 244866 445938 245102 446174
rect 244546 445618 244782 445854
rect 244866 445618 245102 445854
rect 244546 405938 244782 406174
rect 244866 405938 245102 406174
rect 244546 405618 244782 405854
rect 244866 405618 245102 405854
rect 244546 365938 244782 366174
rect 244866 365938 245102 366174
rect 244546 365618 244782 365854
rect 244866 365618 245102 365854
rect 244546 325938 244782 326174
rect 244866 325938 245102 326174
rect 244546 325618 244782 325854
rect 244866 325618 245102 325854
rect 244546 285938 244782 286174
rect 244866 285938 245102 286174
rect 244546 285618 244782 285854
rect 244866 285618 245102 285854
rect 244546 245938 244782 246174
rect 244866 245938 245102 246174
rect 244546 245618 244782 245854
rect 244866 245618 245102 245854
rect 244546 205938 244782 206174
rect 244866 205938 245102 206174
rect 244546 205618 244782 205854
rect 244866 205618 245102 205854
rect 244546 165938 244782 166174
rect 244866 165938 245102 166174
rect 244546 165618 244782 165854
rect 244866 165618 245102 165854
rect 244546 125938 244782 126174
rect 244866 125938 245102 126174
rect 244546 125618 244782 125854
rect 244866 125618 245102 125854
rect 244546 85938 244782 86174
rect 244866 85938 245102 86174
rect 244546 85618 244782 85854
rect 244866 85618 245102 85854
rect 244546 45938 244782 46174
rect 244866 45938 245102 46174
rect 244546 45618 244782 45854
rect 244866 45618 245102 45854
rect 244546 5938 244782 6174
rect 244866 5938 245102 6174
rect 244546 5618 244782 5854
rect 244866 5618 245102 5854
rect 244546 -2502 244782 -2266
rect 244866 -2502 245102 -2266
rect 244546 -2822 244782 -2586
rect 244866 -2822 245102 -2586
rect 248266 689658 248502 689894
rect 248586 689658 248822 689894
rect 248266 689338 248502 689574
rect 248586 689338 248822 689574
rect 248266 649658 248502 649894
rect 248586 649658 248822 649894
rect 248266 649338 248502 649574
rect 248586 649338 248822 649574
rect 248266 609658 248502 609894
rect 248586 609658 248822 609894
rect 248266 609338 248502 609574
rect 248586 609338 248822 609574
rect 248266 569658 248502 569894
rect 248586 569658 248822 569894
rect 248266 569338 248502 569574
rect 248586 569338 248822 569574
rect 248266 529658 248502 529894
rect 248586 529658 248822 529894
rect 248266 529338 248502 529574
rect 248586 529338 248822 529574
rect 248266 489658 248502 489894
rect 248586 489658 248822 489894
rect 248266 489338 248502 489574
rect 248586 489338 248822 489574
rect 248266 449658 248502 449894
rect 248586 449658 248822 449894
rect 248266 449338 248502 449574
rect 248586 449338 248822 449574
rect 248266 409658 248502 409894
rect 248586 409658 248822 409894
rect 248266 409338 248502 409574
rect 248586 409338 248822 409574
rect 248266 369658 248502 369894
rect 248586 369658 248822 369894
rect 248266 369338 248502 369574
rect 248586 369338 248822 369574
rect 248266 329658 248502 329894
rect 248586 329658 248822 329894
rect 248266 329338 248502 329574
rect 248586 329338 248822 329574
rect 248266 289658 248502 289894
rect 248586 289658 248822 289894
rect 248266 289338 248502 289574
rect 248586 289338 248822 289574
rect 248266 249658 248502 249894
rect 248586 249658 248822 249894
rect 248266 249338 248502 249574
rect 248586 249338 248822 249574
rect 248266 209658 248502 209894
rect 248586 209658 248822 209894
rect 248266 209338 248502 209574
rect 248586 209338 248822 209574
rect 248266 169658 248502 169894
rect 248586 169658 248822 169894
rect 248266 169338 248502 169574
rect 248586 169338 248822 169574
rect 248266 129658 248502 129894
rect 248586 129658 248822 129894
rect 248266 129338 248502 129574
rect 248586 129338 248822 129574
rect 248266 89658 248502 89894
rect 248586 89658 248822 89894
rect 248266 89338 248502 89574
rect 248586 89338 248822 89574
rect 248266 49658 248502 49894
rect 248586 49658 248822 49894
rect 248266 49338 248502 49574
rect 248586 49338 248822 49574
rect 248266 9658 248502 9894
rect 248586 9658 248822 9894
rect 248266 9338 248502 9574
rect 248586 9338 248822 9574
rect 248266 -4422 248502 -4186
rect 248586 -4422 248822 -4186
rect 248266 -4742 248502 -4506
rect 248586 -4742 248822 -4506
rect 271986 711322 272222 711558
rect 272306 711322 272542 711558
rect 271986 711002 272222 711238
rect 272306 711002 272542 711238
rect 268266 709402 268502 709638
rect 268586 709402 268822 709638
rect 268266 709082 268502 709318
rect 268586 709082 268822 709318
rect 264546 707482 264782 707718
rect 264866 707482 265102 707718
rect 264546 707162 264782 707398
rect 264866 707162 265102 707398
rect 251986 693378 252222 693614
rect 252306 693378 252542 693614
rect 251986 693058 252222 693294
rect 252306 693058 252542 693294
rect 251986 653378 252222 653614
rect 252306 653378 252542 653614
rect 251986 653058 252222 653294
rect 252306 653058 252542 653294
rect 251986 613378 252222 613614
rect 252306 613378 252542 613614
rect 251986 613058 252222 613294
rect 252306 613058 252542 613294
rect 251986 573378 252222 573614
rect 252306 573378 252542 573614
rect 251986 573058 252222 573294
rect 252306 573058 252542 573294
rect 251986 533378 252222 533614
rect 252306 533378 252542 533614
rect 251986 533058 252222 533294
rect 252306 533058 252542 533294
rect 251986 493378 252222 493614
rect 252306 493378 252542 493614
rect 251986 493058 252222 493294
rect 252306 493058 252542 493294
rect 251986 453378 252222 453614
rect 252306 453378 252542 453614
rect 251986 453058 252222 453294
rect 252306 453058 252542 453294
rect 251986 413378 252222 413614
rect 252306 413378 252542 413614
rect 251986 413058 252222 413294
rect 252306 413058 252542 413294
rect 251986 373378 252222 373614
rect 252306 373378 252542 373614
rect 251986 373058 252222 373294
rect 252306 373058 252542 373294
rect 251986 333378 252222 333614
rect 252306 333378 252542 333614
rect 251986 333058 252222 333294
rect 252306 333058 252542 333294
rect 251986 293378 252222 293614
rect 252306 293378 252542 293614
rect 251986 293058 252222 293294
rect 252306 293058 252542 293294
rect 251986 253378 252222 253614
rect 252306 253378 252542 253614
rect 251986 253058 252222 253294
rect 252306 253058 252542 253294
rect 251986 213378 252222 213614
rect 252306 213378 252542 213614
rect 251986 213058 252222 213294
rect 252306 213058 252542 213294
rect 251986 173378 252222 173614
rect 252306 173378 252542 173614
rect 251986 173058 252222 173294
rect 252306 173058 252542 173294
rect 251986 133378 252222 133614
rect 252306 133378 252542 133614
rect 251986 133058 252222 133294
rect 252306 133058 252542 133294
rect 251986 93378 252222 93614
rect 252306 93378 252542 93614
rect 251986 93058 252222 93294
rect 252306 93058 252542 93294
rect 251986 53378 252222 53614
rect 252306 53378 252542 53614
rect 251986 53058 252222 53294
rect 252306 53058 252542 53294
rect 251986 13378 252222 13614
rect 252306 13378 252542 13614
rect 251986 13058 252222 13294
rect 252306 13058 252542 13294
rect 231986 -7302 232222 -7066
rect 232306 -7302 232542 -7066
rect 231986 -7622 232222 -7386
rect 232306 -7622 232542 -7386
rect 260826 705562 261062 705798
rect 261146 705562 261382 705798
rect 260826 705242 261062 705478
rect 261146 705242 261382 705478
rect 260826 662218 261062 662454
rect 261146 662218 261382 662454
rect 260826 661898 261062 662134
rect 261146 661898 261382 662134
rect 260826 622218 261062 622454
rect 261146 622218 261382 622454
rect 260826 621898 261062 622134
rect 261146 621898 261382 622134
rect 260826 582218 261062 582454
rect 261146 582218 261382 582454
rect 260826 581898 261062 582134
rect 261146 581898 261382 582134
rect 260826 542218 261062 542454
rect 261146 542218 261382 542454
rect 260826 541898 261062 542134
rect 261146 541898 261382 542134
rect 260826 502218 261062 502454
rect 261146 502218 261382 502454
rect 260826 501898 261062 502134
rect 261146 501898 261382 502134
rect 260826 462218 261062 462454
rect 261146 462218 261382 462454
rect 260826 461898 261062 462134
rect 261146 461898 261382 462134
rect 260826 422218 261062 422454
rect 261146 422218 261382 422454
rect 260826 421898 261062 422134
rect 261146 421898 261382 422134
rect 260826 382218 261062 382454
rect 261146 382218 261382 382454
rect 260826 381898 261062 382134
rect 261146 381898 261382 382134
rect 260826 342218 261062 342454
rect 261146 342218 261382 342454
rect 260826 341898 261062 342134
rect 261146 341898 261382 342134
rect 260826 302218 261382 302454
rect 260826 301898 261382 302134
rect 260826 262218 261382 262454
rect 260826 261898 261382 262134
rect 260826 222218 261382 222454
rect 260826 221898 261382 222134
rect 260826 182218 261382 182454
rect 260826 181898 261382 182134
rect 260826 142218 261382 142454
rect 260826 141898 261382 142134
rect 260826 102218 261062 102454
rect 261146 102218 261382 102454
rect 260826 101898 261062 102134
rect 261146 101898 261382 102134
rect 260826 62218 261062 62454
rect 261146 62218 261382 62454
rect 260826 61898 261062 62134
rect 261146 61898 261382 62134
rect 260826 22218 261062 22454
rect 261146 22218 261382 22454
rect 260826 21898 261062 22134
rect 261146 21898 261382 22134
rect 260826 -1542 261062 -1306
rect 261146 -1542 261382 -1306
rect 260826 -1862 261062 -1626
rect 261146 -1862 261382 -1626
rect 264546 665938 264782 666174
rect 264866 665938 265102 666174
rect 264546 665618 264782 665854
rect 264866 665618 265102 665854
rect 264546 625938 264782 626174
rect 264866 625938 265102 626174
rect 264546 625618 264782 625854
rect 264866 625618 265102 625854
rect 264546 585938 264782 586174
rect 264866 585938 265102 586174
rect 264546 585618 264782 585854
rect 264866 585618 265102 585854
rect 264546 545938 264782 546174
rect 264866 545938 265102 546174
rect 264546 545618 264782 545854
rect 264866 545618 265102 545854
rect 264546 505938 264782 506174
rect 264866 505938 265102 506174
rect 264546 505618 264782 505854
rect 264866 505618 265102 505854
rect 264546 465938 264782 466174
rect 264866 465938 265102 466174
rect 264546 465618 264782 465854
rect 264866 465618 265102 465854
rect 264546 425938 264782 426174
rect 264866 425938 265102 426174
rect 264546 425618 264782 425854
rect 264866 425618 265102 425854
rect 264546 385938 264782 386174
rect 264866 385938 265102 386174
rect 264546 385618 264782 385854
rect 264866 385618 265102 385854
rect 264546 345938 264782 346174
rect 264866 345938 265102 346174
rect 264546 345618 264782 345854
rect 264866 345618 265102 345854
rect 264546 305938 264782 306174
rect 264866 305938 265102 306174
rect 264546 305618 264782 305854
rect 264866 305618 265102 305854
rect 264546 265938 264782 266174
rect 264866 265938 265102 266174
rect 264546 265618 264782 265854
rect 264866 265618 265102 265854
rect 264546 225938 264782 226174
rect 264866 225938 265102 226174
rect 264546 225618 264782 225854
rect 264866 225618 265102 225854
rect 264546 185938 264782 186174
rect 264866 185938 265102 186174
rect 264546 185618 264782 185854
rect 264866 185618 265102 185854
rect 264546 145938 264782 146174
rect 264866 145938 265102 146174
rect 264546 145618 264782 145854
rect 264866 145618 265102 145854
rect 264546 105938 264782 106174
rect 264866 105938 265102 106174
rect 264546 105618 264782 105854
rect 264866 105618 265102 105854
rect 264546 65938 264782 66174
rect 264866 65938 265102 66174
rect 264546 65618 264782 65854
rect 264866 65618 265102 65854
rect 264546 25938 264782 26174
rect 264866 25938 265102 26174
rect 264546 25618 264782 25854
rect 264866 25618 265102 25854
rect 264546 -3462 264782 -3226
rect 264866 -3462 265102 -3226
rect 264546 -3782 264782 -3546
rect 264866 -3782 265102 -3546
rect 268266 669658 268502 669894
rect 268586 669658 268822 669894
rect 268266 669338 268502 669574
rect 268586 669338 268822 669574
rect 268266 629658 268502 629894
rect 268586 629658 268822 629894
rect 268266 629338 268502 629574
rect 268586 629338 268822 629574
rect 268266 589658 268502 589894
rect 268586 589658 268822 589894
rect 268266 589338 268502 589574
rect 268586 589338 268822 589574
rect 268266 549658 268502 549894
rect 268586 549658 268822 549894
rect 268266 549338 268502 549574
rect 268586 549338 268822 549574
rect 268266 509658 268502 509894
rect 268586 509658 268822 509894
rect 268266 509338 268502 509574
rect 268586 509338 268822 509574
rect 268266 469658 268502 469894
rect 268586 469658 268822 469894
rect 268266 469338 268502 469574
rect 268586 469338 268822 469574
rect 268266 429658 268502 429894
rect 268586 429658 268822 429894
rect 268266 429338 268502 429574
rect 268586 429338 268822 429574
rect 268266 389658 268502 389894
rect 268586 389658 268822 389894
rect 268266 389338 268502 389574
rect 268586 389338 268822 389574
rect 268266 349658 268502 349894
rect 268586 349658 268822 349894
rect 268266 349338 268502 349574
rect 268586 349338 268822 349574
rect 268266 309658 268502 309894
rect 268586 309658 268822 309894
rect 268266 309338 268502 309574
rect 268586 309338 268822 309574
rect 268266 269658 268502 269894
rect 268586 269658 268822 269894
rect 268266 269338 268502 269574
rect 268586 269338 268822 269574
rect 268266 229658 268502 229894
rect 268586 229658 268822 229894
rect 268266 229338 268502 229574
rect 268586 229338 268822 229574
rect 268266 189658 268502 189894
rect 268586 189658 268822 189894
rect 268266 189338 268502 189574
rect 268586 189338 268822 189574
rect 268266 149658 268502 149894
rect 268586 149658 268822 149894
rect 268266 149338 268502 149574
rect 268586 149338 268822 149574
rect 268266 109658 268502 109894
rect 268586 109658 268822 109894
rect 268266 109338 268502 109574
rect 268586 109338 268822 109574
rect 268266 69658 268502 69894
rect 268586 69658 268822 69894
rect 268266 69338 268502 69574
rect 268586 69338 268822 69574
rect 268266 29658 268502 29894
rect 268586 29658 268822 29894
rect 268266 29338 268502 29574
rect 268586 29338 268822 29574
rect 268266 -5382 268502 -5146
rect 268586 -5382 268822 -5146
rect 268266 -5702 268502 -5466
rect 268586 -5702 268822 -5466
rect 291986 710362 292222 710598
rect 292306 710362 292542 710598
rect 291986 710042 292222 710278
rect 292306 710042 292542 710278
rect 288266 708442 288502 708678
rect 288586 708442 288822 708678
rect 288266 708122 288502 708358
rect 288586 708122 288822 708358
rect 284546 706522 284782 706758
rect 284866 706522 285102 706758
rect 284546 706202 284782 706438
rect 284866 706202 285102 706438
rect 271986 673378 272222 673614
rect 272306 673378 272542 673614
rect 271986 673058 272222 673294
rect 272306 673058 272542 673294
rect 271986 633378 272222 633614
rect 272306 633378 272542 633614
rect 271986 633058 272222 633294
rect 272306 633058 272542 633294
rect 271986 593378 272222 593614
rect 272306 593378 272542 593614
rect 271986 593058 272222 593294
rect 272306 593058 272542 593294
rect 271986 553378 272222 553614
rect 272306 553378 272542 553614
rect 271986 553058 272222 553294
rect 272306 553058 272542 553294
rect 271986 513378 272222 513614
rect 272306 513378 272542 513614
rect 271986 513058 272222 513294
rect 272306 513058 272542 513294
rect 271986 473378 272222 473614
rect 272306 473378 272542 473614
rect 271986 473058 272222 473294
rect 272306 473058 272542 473294
rect 271986 433378 272222 433614
rect 272306 433378 272542 433614
rect 271986 433058 272222 433294
rect 272306 433058 272542 433294
rect 271986 393378 272222 393614
rect 272306 393378 272542 393614
rect 271986 393058 272222 393294
rect 272306 393058 272542 393294
rect 271986 353378 272222 353614
rect 272306 353378 272542 353614
rect 271986 353058 272222 353294
rect 272306 353058 272542 353294
rect 280826 704602 281062 704838
rect 281146 704602 281382 704838
rect 280826 704282 281062 704518
rect 281146 704282 281382 704518
rect 280826 682218 281062 682454
rect 281146 682218 281382 682454
rect 280826 681898 281062 682134
rect 281146 681898 281382 682134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 602218 281062 602454
rect 281146 602218 281382 602454
rect 280826 601898 281062 602134
rect 281146 601898 281382 602134
rect 280826 562218 281062 562454
rect 281146 562218 281382 562454
rect 280826 561898 281062 562134
rect 281146 561898 281382 562134
rect 280826 522218 281062 522454
rect 281146 522218 281382 522454
rect 280826 521898 281062 522134
rect 281146 521898 281382 522134
rect 280826 482218 281062 482454
rect 281146 482218 281382 482454
rect 280826 481898 281062 482134
rect 281146 481898 281382 482134
rect 280826 442218 281062 442454
rect 281146 442218 281382 442454
rect 280826 441898 281062 442134
rect 281146 441898 281382 442134
rect 280826 402218 281062 402454
rect 281146 402218 281382 402454
rect 280826 401898 281062 402134
rect 281146 401898 281382 402134
rect 280826 362218 281062 362454
rect 281146 362218 281382 362454
rect 280826 361898 281062 362134
rect 281146 361898 281382 362134
rect 280826 322218 281062 322454
rect 281146 322218 281382 322454
rect 280826 321898 281062 322134
rect 281146 321898 281382 322134
rect 271986 313378 272222 313614
rect 272306 313378 272542 313614
rect 271986 313058 272222 313294
rect 272306 313058 272542 313294
rect 271986 273378 272222 273614
rect 272306 273378 272542 273614
rect 271986 273058 272222 273294
rect 272306 273058 272542 273294
rect 271986 233378 272222 233614
rect 272306 233378 272542 233614
rect 271986 233058 272222 233294
rect 272306 233058 272542 233294
rect 271986 193378 272222 193614
rect 272306 193378 272542 193614
rect 271986 193058 272222 193294
rect 272306 193058 272542 193294
rect 271986 153378 272222 153614
rect 272306 153378 272542 153614
rect 271986 153058 272222 153294
rect 272306 153058 272542 153294
rect 271986 113378 272222 113614
rect 272306 113378 272542 113614
rect 271986 113058 272222 113294
rect 272306 113058 272542 113294
rect 271986 73378 272222 73614
rect 272306 73378 272542 73614
rect 271986 73058 272222 73294
rect 272306 73058 272542 73294
rect 271986 33378 272222 33614
rect 272306 33378 272542 33614
rect 271986 33058 272222 33294
rect 272306 33058 272542 33294
rect 251986 -6342 252222 -6106
rect 252306 -6342 252542 -6106
rect 251986 -6662 252222 -6426
rect 252306 -6662 252542 -6426
rect 284546 685938 284782 686174
rect 284866 685938 285102 686174
rect 284546 685618 284782 685854
rect 284866 685618 285102 685854
rect 284546 645938 284782 646174
rect 284866 645938 285102 646174
rect 284546 645618 284782 645854
rect 284866 645618 285102 645854
rect 284546 605938 284782 606174
rect 284866 605938 285102 606174
rect 284546 605618 284782 605854
rect 284866 605618 285102 605854
rect 284546 565938 284782 566174
rect 284866 565938 285102 566174
rect 284546 565618 284782 565854
rect 284866 565618 285102 565854
rect 284546 525938 284782 526174
rect 284866 525938 285102 526174
rect 284546 525618 284782 525854
rect 284866 525618 285102 525854
rect 284546 485938 284782 486174
rect 284866 485938 285102 486174
rect 284546 485618 284782 485854
rect 284866 485618 285102 485854
rect 284546 445938 284782 446174
rect 284866 445938 285102 446174
rect 284546 445618 284782 445854
rect 284866 445618 285102 445854
rect 284546 405938 284782 406174
rect 284866 405938 285102 406174
rect 284546 405618 284782 405854
rect 284866 405618 285102 405854
rect 284546 365938 284782 366174
rect 284866 365938 285102 366174
rect 284546 365618 284782 365854
rect 284866 365618 285102 365854
rect 284546 325938 284782 326174
rect 284866 325938 285102 326174
rect 284546 325618 284782 325854
rect 284866 325618 285102 325854
rect 280826 282218 281382 282454
rect 280826 281898 281382 282134
rect 280826 242218 281382 242454
rect 280826 241898 281382 242134
rect 280826 202218 281382 202454
rect 280826 201898 281382 202134
rect 280826 162218 281382 162454
rect 280826 161898 281382 162134
rect 280826 122218 281062 122454
rect 281146 122218 281382 122454
rect 280826 121898 281062 122134
rect 281146 121898 281382 122134
rect 280826 82218 281062 82454
rect 281146 82218 281382 82454
rect 280826 81898 281062 82134
rect 281146 81898 281382 82134
rect 280826 42218 281062 42454
rect 281146 42218 281382 42454
rect 280826 41898 281062 42134
rect 281146 41898 281382 42134
rect 284546 285938 284782 286174
rect 284866 285938 285102 286174
rect 284546 285618 284782 285854
rect 284866 285618 285102 285854
rect 284546 245938 284782 246174
rect 284866 245938 285102 246174
rect 284546 245618 284782 245854
rect 284866 245618 285102 245854
rect 284546 205938 284782 206174
rect 284866 205938 285102 206174
rect 284546 205618 284782 205854
rect 284866 205618 285102 205854
rect 284546 165938 284782 166174
rect 284866 165938 285102 166174
rect 284546 165618 284782 165854
rect 284866 165618 285102 165854
rect 284546 125938 284782 126174
rect 284866 125938 285102 126174
rect 284546 125618 284782 125854
rect 284866 125618 285102 125854
rect 284546 85938 284782 86174
rect 284866 85938 285102 86174
rect 284546 85618 284782 85854
rect 284866 85618 285102 85854
rect 284546 45938 284782 46174
rect 284866 45938 285102 46174
rect 284546 45618 284782 45854
rect 284866 45618 285102 45854
rect 284546 5938 284782 6174
rect 284866 5938 285102 6174
rect 284546 5618 284782 5854
rect 284866 5618 285102 5854
rect 280826 2218 281062 2454
rect 281146 2218 281382 2454
rect 280826 1898 281062 2134
rect 281146 1898 281382 2134
rect 280826 -582 281062 -346
rect 281146 -582 281382 -346
rect 280826 -902 281062 -666
rect 281146 -902 281382 -666
rect 284546 -2502 284782 -2266
rect 284866 -2502 285102 -2266
rect 284546 -2822 284782 -2586
rect 284866 -2822 285102 -2586
rect 288266 689658 288502 689894
rect 288586 689658 288822 689894
rect 288266 689338 288502 689574
rect 288586 689338 288822 689574
rect 288266 649658 288502 649894
rect 288586 649658 288822 649894
rect 288266 649338 288502 649574
rect 288586 649338 288822 649574
rect 288266 609658 288502 609894
rect 288586 609658 288822 609894
rect 288266 609338 288502 609574
rect 288586 609338 288822 609574
rect 288266 569658 288502 569894
rect 288586 569658 288822 569894
rect 288266 569338 288502 569574
rect 288586 569338 288822 569574
rect 288266 529658 288502 529894
rect 288586 529658 288822 529894
rect 288266 529338 288502 529574
rect 288586 529338 288822 529574
rect 288266 489658 288502 489894
rect 288586 489658 288822 489894
rect 288266 489338 288502 489574
rect 288586 489338 288822 489574
rect 288266 449658 288502 449894
rect 288586 449658 288822 449894
rect 288266 449338 288502 449574
rect 288586 449338 288822 449574
rect 288266 409658 288502 409894
rect 288586 409658 288822 409894
rect 288266 409338 288502 409574
rect 288586 409338 288822 409574
rect 288266 369658 288502 369894
rect 288586 369658 288822 369894
rect 288266 369338 288502 369574
rect 288586 369338 288822 369574
rect 288266 329658 288502 329894
rect 288586 329658 288822 329894
rect 288266 329338 288502 329574
rect 288586 329338 288822 329574
rect 288266 289658 288502 289894
rect 288586 289658 288822 289894
rect 288266 289338 288502 289574
rect 288586 289338 288822 289574
rect 288266 249658 288502 249894
rect 288586 249658 288822 249894
rect 288266 249338 288502 249574
rect 288586 249338 288822 249574
rect 288266 209658 288502 209894
rect 288586 209658 288822 209894
rect 288266 209338 288502 209574
rect 288586 209338 288822 209574
rect 288266 169658 288502 169894
rect 288586 169658 288822 169894
rect 288266 169338 288502 169574
rect 288586 169338 288822 169574
rect 288266 129658 288502 129894
rect 288586 129658 288822 129894
rect 288266 129338 288502 129574
rect 288586 129338 288822 129574
rect 288266 89658 288502 89894
rect 288586 89658 288822 89894
rect 288266 89338 288502 89574
rect 288586 89338 288822 89574
rect 288266 49658 288502 49894
rect 288586 49658 288822 49894
rect 288266 49338 288502 49574
rect 288586 49338 288822 49574
rect 288266 9658 288502 9894
rect 288586 9658 288822 9894
rect 288266 9338 288502 9574
rect 288586 9338 288822 9574
rect 288266 -4422 288502 -4186
rect 288586 -4422 288822 -4186
rect 288266 -4742 288502 -4506
rect 288586 -4742 288822 -4506
rect 311986 711322 312222 711558
rect 312306 711322 312542 711558
rect 311986 711002 312222 711238
rect 312306 711002 312542 711238
rect 308266 709402 308502 709638
rect 308586 709402 308822 709638
rect 308266 709082 308502 709318
rect 308586 709082 308822 709318
rect 304546 707482 304782 707718
rect 304866 707482 305102 707718
rect 304546 707162 304782 707398
rect 304866 707162 305102 707398
rect 291986 693378 292222 693614
rect 292306 693378 292542 693614
rect 291986 693058 292222 693294
rect 292306 693058 292542 693294
rect 291986 653378 292222 653614
rect 292306 653378 292542 653614
rect 291986 653058 292222 653294
rect 292306 653058 292542 653294
rect 291986 613378 292222 613614
rect 292306 613378 292542 613614
rect 291986 613058 292222 613294
rect 292306 613058 292542 613294
rect 291986 573378 292222 573614
rect 292306 573378 292542 573614
rect 291986 573058 292222 573294
rect 292306 573058 292542 573294
rect 291986 533378 292222 533614
rect 292306 533378 292542 533614
rect 291986 533058 292222 533294
rect 292306 533058 292542 533294
rect 291986 493378 292222 493614
rect 292306 493378 292542 493614
rect 291986 493058 292222 493294
rect 292306 493058 292542 493294
rect 291986 453378 292222 453614
rect 292306 453378 292542 453614
rect 291986 453058 292222 453294
rect 292306 453058 292542 453294
rect 291986 413378 292222 413614
rect 292306 413378 292542 413614
rect 291986 413058 292222 413294
rect 292306 413058 292542 413294
rect 291986 373378 292222 373614
rect 292306 373378 292542 373614
rect 291986 373058 292222 373294
rect 292306 373058 292542 373294
rect 291986 333378 292222 333614
rect 292306 333378 292542 333614
rect 291986 333058 292222 333294
rect 292306 333058 292542 333294
rect 300826 705562 301062 705798
rect 301146 705562 301382 705798
rect 300826 705242 301062 705478
rect 301146 705242 301382 705478
rect 300826 662218 301062 662454
rect 301146 662218 301382 662454
rect 300826 661898 301062 662134
rect 301146 661898 301382 662134
rect 300826 622218 301062 622454
rect 301146 622218 301382 622454
rect 300826 621898 301062 622134
rect 301146 621898 301382 622134
rect 300826 582218 301062 582454
rect 301146 582218 301382 582454
rect 300826 581898 301062 582134
rect 301146 581898 301382 582134
rect 300826 542218 301062 542454
rect 301146 542218 301382 542454
rect 300826 541898 301062 542134
rect 301146 541898 301382 542134
rect 300826 502218 301062 502454
rect 301146 502218 301382 502454
rect 300826 501898 301062 502134
rect 301146 501898 301382 502134
rect 300826 462218 301062 462454
rect 301146 462218 301382 462454
rect 300826 461898 301062 462134
rect 301146 461898 301382 462134
rect 300826 422218 301062 422454
rect 301146 422218 301382 422454
rect 300826 421898 301062 422134
rect 301146 421898 301382 422134
rect 300826 382218 301062 382454
rect 301146 382218 301382 382454
rect 300826 381898 301062 382134
rect 301146 381898 301382 382134
rect 300826 342218 301062 342454
rect 301146 342218 301382 342454
rect 300826 341898 301062 342134
rect 301146 341898 301382 342134
rect 291986 293378 292222 293614
rect 292306 293378 292542 293614
rect 291986 293058 292222 293294
rect 292306 293058 292542 293294
rect 291986 253378 292222 253614
rect 292306 253378 292542 253614
rect 291986 253058 292222 253294
rect 292306 253058 292542 253294
rect 291986 213378 292222 213614
rect 292306 213378 292542 213614
rect 291986 213058 292222 213294
rect 292306 213058 292542 213294
rect 291986 173378 292222 173614
rect 292306 173378 292542 173614
rect 291986 173058 292222 173294
rect 292306 173058 292542 173294
rect 291986 133378 292222 133614
rect 292306 133378 292542 133614
rect 291986 133058 292222 133294
rect 292306 133058 292542 133294
rect 291986 93378 292222 93614
rect 292306 93378 292542 93614
rect 291986 93058 292222 93294
rect 292306 93058 292542 93294
rect 291986 53378 292222 53614
rect 292306 53378 292542 53614
rect 291986 53058 292222 53294
rect 292306 53058 292542 53294
rect 291986 13378 292222 13614
rect 292306 13378 292542 13614
rect 291986 13058 292222 13294
rect 292306 13058 292542 13294
rect 271986 -7302 272222 -7066
rect 272306 -7302 272542 -7066
rect 271986 -7622 272222 -7386
rect 272306 -7622 272542 -7386
rect 304546 665938 304782 666174
rect 304866 665938 305102 666174
rect 304546 665618 304782 665854
rect 304866 665618 305102 665854
rect 304546 625938 304782 626174
rect 304866 625938 305102 626174
rect 304546 625618 304782 625854
rect 304866 625618 305102 625854
rect 304546 585938 304782 586174
rect 304866 585938 305102 586174
rect 304546 585618 304782 585854
rect 304866 585618 305102 585854
rect 304546 545938 304782 546174
rect 304866 545938 305102 546174
rect 304546 545618 304782 545854
rect 304866 545618 305102 545854
rect 304546 505938 304782 506174
rect 304866 505938 305102 506174
rect 304546 505618 304782 505854
rect 304866 505618 305102 505854
rect 304546 465938 304782 466174
rect 304866 465938 305102 466174
rect 304546 465618 304782 465854
rect 304866 465618 305102 465854
rect 304546 425938 304782 426174
rect 304866 425938 305102 426174
rect 304546 425618 304782 425854
rect 304866 425618 305102 425854
rect 304546 385938 304782 386174
rect 304866 385938 305102 386174
rect 304546 385618 304782 385854
rect 304866 385618 305102 385854
rect 304546 345938 304782 346174
rect 304866 345938 305102 346174
rect 304546 345618 304782 345854
rect 304866 345618 305102 345854
rect 300826 302218 301382 302454
rect 300826 301898 301382 302134
rect 300826 262218 301382 262454
rect 300826 261898 301382 262134
rect 300826 222218 301382 222454
rect 300826 221898 301382 222134
rect 300826 182218 301382 182454
rect 300826 181898 301382 182134
rect 300826 142218 301382 142454
rect 300826 141898 301382 142134
rect 300826 102218 301062 102454
rect 301146 102218 301382 102454
rect 300826 101898 301062 102134
rect 301146 101898 301382 102134
rect 300826 62218 301062 62454
rect 301146 62218 301382 62454
rect 300826 61898 301062 62134
rect 301146 61898 301382 62134
rect 300826 22218 301062 22454
rect 301146 22218 301382 22454
rect 300826 21898 301062 22134
rect 301146 21898 301382 22134
rect 304546 305938 304782 306174
rect 304866 305938 305102 306174
rect 304546 305618 304782 305854
rect 304866 305618 305102 305854
rect 304546 265938 304782 266174
rect 304866 265938 305102 266174
rect 304546 265618 304782 265854
rect 304866 265618 305102 265854
rect 304546 225938 304782 226174
rect 304866 225938 305102 226174
rect 304546 225618 304782 225854
rect 304866 225618 305102 225854
rect 304546 185938 304782 186174
rect 304866 185938 305102 186174
rect 304546 185618 304782 185854
rect 304866 185618 305102 185854
rect 304546 145938 304782 146174
rect 304866 145938 305102 146174
rect 304546 145618 304782 145854
rect 304866 145618 305102 145854
rect 304546 105938 304782 106174
rect 304866 105938 305102 106174
rect 304546 105618 304782 105854
rect 304866 105618 305102 105854
rect 304546 65938 304782 66174
rect 304866 65938 305102 66174
rect 304546 65618 304782 65854
rect 304866 65618 305102 65854
rect 304546 25938 304782 26174
rect 304866 25938 305102 26174
rect 304546 25618 304782 25854
rect 304866 25618 305102 25854
rect 300826 -1542 301062 -1306
rect 301146 -1542 301382 -1306
rect 300826 -1862 301062 -1626
rect 301146 -1862 301382 -1626
rect 304546 -3462 304782 -3226
rect 304866 -3462 305102 -3226
rect 304546 -3782 304782 -3546
rect 304866 -3782 305102 -3546
rect 308266 669658 308502 669894
rect 308586 669658 308822 669894
rect 308266 669338 308502 669574
rect 308586 669338 308822 669574
rect 308266 629658 308502 629894
rect 308586 629658 308822 629894
rect 308266 629338 308502 629574
rect 308586 629338 308822 629574
rect 308266 589658 308502 589894
rect 308586 589658 308822 589894
rect 308266 589338 308502 589574
rect 308586 589338 308822 589574
rect 308266 549658 308502 549894
rect 308586 549658 308822 549894
rect 308266 549338 308502 549574
rect 308586 549338 308822 549574
rect 308266 509658 308502 509894
rect 308586 509658 308822 509894
rect 308266 509338 308502 509574
rect 308586 509338 308822 509574
rect 308266 469658 308502 469894
rect 308586 469658 308822 469894
rect 308266 469338 308502 469574
rect 308586 469338 308822 469574
rect 308266 429658 308502 429894
rect 308586 429658 308822 429894
rect 308266 429338 308502 429574
rect 308586 429338 308822 429574
rect 308266 389658 308502 389894
rect 308586 389658 308822 389894
rect 308266 389338 308502 389574
rect 308586 389338 308822 389574
rect 308266 349658 308502 349894
rect 308586 349658 308822 349894
rect 308266 349338 308502 349574
rect 308586 349338 308822 349574
rect 308266 309658 308502 309894
rect 308586 309658 308822 309894
rect 308266 309338 308502 309574
rect 308586 309338 308822 309574
rect 308266 269658 308502 269894
rect 308586 269658 308822 269894
rect 308266 269338 308502 269574
rect 308586 269338 308822 269574
rect 308266 229658 308502 229894
rect 308586 229658 308822 229894
rect 308266 229338 308502 229574
rect 308586 229338 308822 229574
rect 308266 189658 308502 189894
rect 308586 189658 308822 189894
rect 308266 189338 308502 189574
rect 308586 189338 308822 189574
rect 308266 149658 308502 149894
rect 308586 149658 308822 149894
rect 308266 149338 308502 149574
rect 308586 149338 308822 149574
rect 308266 109658 308502 109894
rect 308586 109658 308822 109894
rect 308266 109338 308502 109574
rect 308586 109338 308822 109574
rect 308266 69658 308502 69894
rect 308586 69658 308822 69894
rect 308266 69338 308502 69574
rect 308586 69338 308822 69574
rect 308266 29658 308502 29894
rect 308586 29658 308822 29894
rect 308266 29338 308502 29574
rect 308586 29338 308822 29574
rect 308266 -5382 308502 -5146
rect 308586 -5382 308822 -5146
rect 308266 -5702 308502 -5466
rect 308586 -5702 308822 -5466
rect 331986 710362 332222 710598
rect 332306 710362 332542 710598
rect 331986 710042 332222 710278
rect 332306 710042 332542 710278
rect 328266 708442 328502 708678
rect 328586 708442 328822 708678
rect 328266 708122 328502 708358
rect 328586 708122 328822 708358
rect 324546 706522 324782 706758
rect 324866 706522 325102 706758
rect 324546 706202 324782 706438
rect 324866 706202 325102 706438
rect 311986 673378 312222 673614
rect 312306 673378 312542 673614
rect 311986 673058 312222 673294
rect 312306 673058 312542 673294
rect 311986 633378 312222 633614
rect 312306 633378 312542 633614
rect 311986 633058 312222 633294
rect 312306 633058 312542 633294
rect 311986 593378 312222 593614
rect 312306 593378 312542 593614
rect 311986 593058 312222 593294
rect 312306 593058 312542 593294
rect 311986 553378 312222 553614
rect 312306 553378 312542 553614
rect 311986 553058 312222 553294
rect 312306 553058 312542 553294
rect 311986 513378 312222 513614
rect 312306 513378 312542 513614
rect 311986 513058 312222 513294
rect 312306 513058 312542 513294
rect 311986 473378 312222 473614
rect 312306 473378 312542 473614
rect 311986 473058 312222 473294
rect 312306 473058 312542 473294
rect 311986 433378 312222 433614
rect 312306 433378 312542 433614
rect 311986 433058 312222 433294
rect 312306 433058 312542 433294
rect 311986 393378 312222 393614
rect 312306 393378 312542 393614
rect 311986 393058 312222 393294
rect 312306 393058 312542 393294
rect 311986 353378 312222 353614
rect 312306 353378 312542 353614
rect 311986 353058 312222 353294
rect 312306 353058 312542 353294
rect 320826 704602 321062 704838
rect 321146 704602 321382 704838
rect 320826 704282 321062 704518
rect 321146 704282 321382 704518
rect 320826 682218 321062 682454
rect 321146 682218 321382 682454
rect 320826 681898 321062 682134
rect 321146 681898 321382 682134
rect 320826 642218 321062 642454
rect 321146 642218 321382 642454
rect 320826 641898 321062 642134
rect 321146 641898 321382 642134
rect 320826 602218 321062 602454
rect 321146 602218 321382 602454
rect 320826 601898 321062 602134
rect 321146 601898 321382 602134
rect 320826 562218 321062 562454
rect 321146 562218 321382 562454
rect 320826 561898 321062 562134
rect 321146 561898 321382 562134
rect 320826 522218 321062 522454
rect 321146 522218 321382 522454
rect 320826 521898 321062 522134
rect 321146 521898 321382 522134
rect 320826 482218 321062 482454
rect 321146 482218 321382 482454
rect 320826 481898 321062 482134
rect 321146 481898 321382 482134
rect 320826 442218 321062 442454
rect 321146 442218 321382 442454
rect 320826 441898 321062 442134
rect 321146 441898 321382 442134
rect 320826 402218 321062 402454
rect 321146 402218 321382 402454
rect 320826 401898 321062 402134
rect 321146 401898 321382 402134
rect 320826 362218 321062 362454
rect 321146 362218 321382 362454
rect 320826 361898 321062 362134
rect 321146 361898 321382 362134
rect 320826 322218 321062 322454
rect 321146 322218 321382 322454
rect 320826 321898 321062 322134
rect 321146 321898 321382 322134
rect 311986 313378 312222 313614
rect 312306 313378 312542 313614
rect 311986 313058 312222 313294
rect 312306 313058 312542 313294
rect 311986 273378 312222 273614
rect 312306 273378 312542 273614
rect 311986 273058 312222 273294
rect 312306 273058 312542 273294
rect 311986 233378 312222 233614
rect 312306 233378 312542 233614
rect 311986 233058 312222 233294
rect 312306 233058 312542 233294
rect 311986 193378 312222 193614
rect 312306 193378 312542 193614
rect 311986 193058 312222 193294
rect 312306 193058 312542 193294
rect 311986 153378 312222 153614
rect 312306 153378 312542 153614
rect 311986 153058 312222 153294
rect 312306 153058 312542 153294
rect 311986 113378 312222 113614
rect 312306 113378 312542 113614
rect 311986 113058 312222 113294
rect 312306 113058 312542 113294
rect 311986 73378 312222 73614
rect 312306 73378 312542 73614
rect 311986 73058 312222 73294
rect 312306 73058 312542 73294
rect 311986 33378 312222 33614
rect 312306 33378 312542 33614
rect 311986 33058 312222 33294
rect 312306 33058 312542 33294
rect 291986 -6342 292222 -6106
rect 292306 -6342 292542 -6106
rect 291986 -6662 292222 -6426
rect 292306 -6662 292542 -6426
rect 320826 282218 321062 282454
rect 321146 282218 321382 282454
rect 320826 281898 321062 282134
rect 321146 281898 321382 282134
rect 320826 242218 321062 242454
rect 321146 242218 321382 242454
rect 320826 241898 321062 242134
rect 321146 241898 321382 242134
rect 320826 202218 321062 202454
rect 321146 202218 321382 202454
rect 320826 201898 321062 202134
rect 321146 201898 321382 202134
rect 320826 162218 321062 162454
rect 321146 162218 321382 162454
rect 320826 161898 321062 162134
rect 321146 161898 321382 162134
rect 320826 122218 321062 122454
rect 321146 122218 321382 122454
rect 320826 121898 321062 122134
rect 321146 121898 321382 122134
rect 320826 82218 321062 82454
rect 321146 82218 321382 82454
rect 320826 81898 321062 82134
rect 321146 81898 321382 82134
rect 320826 42218 321062 42454
rect 321146 42218 321382 42454
rect 320826 41898 321062 42134
rect 321146 41898 321382 42134
rect 320826 2218 321062 2454
rect 321146 2218 321382 2454
rect 320826 1898 321062 2134
rect 321146 1898 321382 2134
rect 320826 -582 321062 -346
rect 321146 -582 321382 -346
rect 320826 -902 321062 -666
rect 321146 -902 321382 -666
rect 324546 685938 324782 686174
rect 324866 685938 325102 686174
rect 324546 685618 324782 685854
rect 324866 685618 325102 685854
rect 324546 645938 324782 646174
rect 324866 645938 325102 646174
rect 324546 645618 324782 645854
rect 324866 645618 325102 645854
rect 324546 605938 324782 606174
rect 324866 605938 325102 606174
rect 324546 605618 324782 605854
rect 324866 605618 325102 605854
rect 324546 565938 324782 566174
rect 324866 565938 325102 566174
rect 324546 565618 324782 565854
rect 324866 565618 325102 565854
rect 324546 525938 324782 526174
rect 324866 525938 325102 526174
rect 324546 525618 324782 525854
rect 324866 525618 325102 525854
rect 324546 485938 324782 486174
rect 324866 485938 325102 486174
rect 324546 485618 324782 485854
rect 324866 485618 325102 485854
rect 324546 445938 324782 446174
rect 324866 445938 325102 446174
rect 324546 445618 324782 445854
rect 324866 445618 325102 445854
rect 324546 405938 324782 406174
rect 324866 405938 325102 406174
rect 324546 405618 324782 405854
rect 324866 405618 325102 405854
rect 324546 365938 324782 366174
rect 324866 365938 325102 366174
rect 324546 365618 324782 365854
rect 324866 365618 325102 365854
rect 324546 325938 324782 326174
rect 324866 325938 325102 326174
rect 324546 325618 324782 325854
rect 324866 325618 325102 325854
rect 324546 285938 324782 286174
rect 324866 285938 325102 286174
rect 324546 285618 324782 285854
rect 324866 285618 325102 285854
rect 324546 245938 324782 246174
rect 324866 245938 325102 246174
rect 324546 245618 324782 245854
rect 324866 245618 325102 245854
rect 324546 205938 324782 206174
rect 324866 205938 325102 206174
rect 324546 205618 324782 205854
rect 324866 205618 325102 205854
rect 324546 165938 324782 166174
rect 324866 165938 325102 166174
rect 324546 165618 324782 165854
rect 324866 165618 325102 165854
rect 324546 125938 324782 126174
rect 324866 125938 325102 126174
rect 324546 125618 324782 125854
rect 324866 125618 325102 125854
rect 324546 85938 324782 86174
rect 324866 85938 325102 86174
rect 324546 85618 324782 85854
rect 324866 85618 325102 85854
rect 324546 45938 324782 46174
rect 324866 45938 325102 46174
rect 324546 45618 324782 45854
rect 324866 45618 325102 45854
rect 324546 5938 324782 6174
rect 324866 5938 325102 6174
rect 324546 5618 324782 5854
rect 324866 5618 325102 5854
rect 324546 -2502 324782 -2266
rect 324866 -2502 325102 -2266
rect 324546 -2822 324782 -2586
rect 324866 -2822 325102 -2586
rect 328266 689658 328502 689894
rect 328586 689658 328822 689894
rect 328266 689338 328502 689574
rect 328586 689338 328822 689574
rect 328266 649658 328502 649894
rect 328586 649658 328822 649894
rect 328266 649338 328502 649574
rect 328586 649338 328822 649574
rect 328266 609658 328502 609894
rect 328586 609658 328822 609894
rect 328266 609338 328502 609574
rect 328586 609338 328822 609574
rect 328266 569658 328502 569894
rect 328586 569658 328822 569894
rect 328266 569338 328502 569574
rect 328586 569338 328822 569574
rect 328266 529658 328502 529894
rect 328586 529658 328822 529894
rect 328266 529338 328502 529574
rect 328586 529338 328822 529574
rect 328266 489658 328502 489894
rect 328586 489658 328822 489894
rect 328266 489338 328502 489574
rect 328586 489338 328822 489574
rect 328266 449658 328502 449894
rect 328586 449658 328822 449894
rect 328266 449338 328502 449574
rect 328586 449338 328822 449574
rect 328266 409658 328502 409894
rect 328586 409658 328822 409894
rect 328266 409338 328502 409574
rect 328586 409338 328822 409574
rect 328266 369658 328502 369894
rect 328586 369658 328822 369894
rect 328266 369338 328502 369574
rect 328586 369338 328822 369574
rect 328266 329658 328502 329894
rect 328586 329658 328822 329894
rect 328266 329338 328502 329574
rect 328586 329338 328822 329574
rect 328266 289658 328502 289894
rect 328586 289658 328822 289894
rect 328266 289338 328502 289574
rect 328586 289338 328822 289574
rect 328266 249658 328502 249894
rect 328586 249658 328822 249894
rect 328266 249338 328502 249574
rect 328586 249338 328822 249574
rect 328266 209658 328502 209894
rect 328586 209658 328822 209894
rect 328266 209338 328502 209574
rect 328586 209338 328822 209574
rect 328266 169658 328502 169894
rect 328586 169658 328822 169894
rect 328266 169338 328502 169574
rect 328586 169338 328822 169574
rect 328266 129658 328502 129894
rect 328586 129658 328822 129894
rect 328266 129338 328502 129574
rect 328586 129338 328822 129574
rect 328266 89658 328502 89894
rect 328586 89658 328822 89894
rect 328266 89338 328502 89574
rect 328586 89338 328822 89574
rect 328266 49658 328502 49894
rect 328586 49658 328822 49894
rect 328266 49338 328502 49574
rect 328586 49338 328822 49574
rect 328266 9658 328502 9894
rect 328586 9658 328822 9894
rect 328266 9338 328502 9574
rect 328586 9338 328822 9574
rect 328266 -4422 328502 -4186
rect 328586 -4422 328822 -4186
rect 328266 -4742 328502 -4506
rect 328586 -4742 328822 -4506
rect 351986 711322 352222 711558
rect 352306 711322 352542 711558
rect 351986 711002 352222 711238
rect 352306 711002 352542 711238
rect 348266 709402 348502 709638
rect 348586 709402 348822 709638
rect 348266 709082 348502 709318
rect 348586 709082 348822 709318
rect 344546 707482 344782 707718
rect 344866 707482 345102 707718
rect 344546 707162 344782 707398
rect 344866 707162 345102 707398
rect 331986 693378 332222 693614
rect 332306 693378 332542 693614
rect 331986 693058 332222 693294
rect 332306 693058 332542 693294
rect 331986 653378 332222 653614
rect 332306 653378 332542 653614
rect 331986 653058 332222 653294
rect 332306 653058 332542 653294
rect 331986 613378 332222 613614
rect 332306 613378 332542 613614
rect 331986 613058 332222 613294
rect 332306 613058 332542 613294
rect 331986 573378 332222 573614
rect 332306 573378 332542 573614
rect 331986 573058 332222 573294
rect 332306 573058 332542 573294
rect 331986 533378 332222 533614
rect 332306 533378 332542 533614
rect 331986 533058 332222 533294
rect 332306 533058 332542 533294
rect 331986 493378 332222 493614
rect 332306 493378 332542 493614
rect 331986 493058 332222 493294
rect 332306 493058 332542 493294
rect 331986 453378 332222 453614
rect 332306 453378 332542 453614
rect 331986 453058 332222 453294
rect 332306 453058 332542 453294
rect 331986 413378 332222 413614
rect 332306 413378 332542 413614
rect 331986 413058 332222 413294
rect 332306 413058 332542 413294
rect 331986 373378 332222 373614
rect 332306 373378 332542 373614
rect 331986 373058 332222 373294
rect 332306 373058 332542 373294
rect 331986 333378 332222 333614
rect 332306 333378 332542 333614
rect 331986 333058 332222 333294
rect 332306 333058 332542 333294
rect 331986 293378 332222 293614
rect 332306 293378 332542 293614
rect 331986 293058 332222 293294
rect 332306 293058 332542 293294
rect 331986 253378 332222 253614
rect 332306 253378 332542 253614
rect 331986 253058 332222 253294
rect 332306 253058 332542 253294
rect 331986 213378 332222 213614
rect 332306 213378 332542 213614
rect 331986 213058 332222 213294
rect 332306 213058 332542 213294
rect 331986 173378 332222 173614
rect 332306 173378 332542 173614
rect 331986 173058 332222 173294
rect 332306 173058 332542 173294
rect 331986 133378 332222 133614
rect 332306 133378 332542 133614
rect 331986 133058 332222 133294
rect 332306 133058 332542 133294
rect 331986 93378 332222 93614
rect 332306 93378 332542 93614
rect 331986 93058 332222 93294
rect 332306 93058 332542 93294
rect 331986 53378 332222 53614
rect 332306 53378 332542 53614
rect 331986 53058 332222 53294
rect 332306 53058 332542 53294
rect 331986 13378 332222 13614
rect 332306 13378 332542 13614
rect 331986 13058 332222 13294
rect 332306 13058 332542 13294
rect 311986 -7302 312222 -7066
rect 312306 -7302 312542 -7066
rect 311986 -7622 312222 -7386
rect 312306 -7622 312542 -7386
rect 340826 705562 341062 705798
rect 341146 705562 341382 705798
rect 340826 705242 341062 705478
rect 341146 705242 341382 705478
rect 340826 662218 341062 662454
rect 341146 662218 341382 662454
rect 340826 661898 341062 662134
rect 341146 661898 341382 662134
rect 340826 622218 341062 622454
rect 341146 622218 341382 622454
rect 340826 621898 341062 622134
rect 341146 621898 341382 622134
rect 340826 582218 341062 582454
rect 341146 582218 341382 582454
rect 340826 581898 341062 582134
rect 341146 581898 341382 582134
rect 340826 542218 341062 542454
rect 341146 542218 341382 542454
rect 340826 541898 341062 542134
rect 341146 541898 341382 542134
rect 340826 502218 341062 502454
rect 341146 502218 341382 502454
rect 340826 501898 341062 502134
rect 341146 501898 341382 502134
rect 340826 462218 341062 462454
rect 341146 462218 341382 462454
rect 340826 461898 341062 462134
rect 341146 461898 341382 462134
rect 340826 422218 341062 422454
rect 341146 422218 341382 422454
rect 340826 421898 341062 422134
rect 341146 421898 341382 422134
rect 340826 382218 341062 382454
rect 341146 382218 341382 382454
rect 340826 381898 341062 382134
rect 341146 381898 341382 382134
rect 340826 342218 341062 342454
rect 341146 342218 341382 342454
rect 340826 341898 341062 342134
rect 341146 341898 341382 342134
rect 340826 302218 341062 302454
rect 341146 302218 341382 302454
rect 340826 301898 341062 302134
rect 341146 301898 341382 302134
rect 340826 262218 341062 262454
rect 341146 262218 341382 262454
rect 340826 261898 341062 262134
rect 341146 261898 341382 262134
rect 340826 222218 341062 222454
rect 341146 222218 341382 222454
rect 340826 221898 341062 222134
rect 341146 221898 341382 222134
rect 340826 182218 341062 182454
rect 341146 182218 341382 182454
rect 340826 181898 341062 182134
rect 341146 181898 341382 182134
rect 340826 142218 341062 142454
rect 341146 142218 341382 142454
rect 340826 141898 341062 142134
rect 341146 141898 341382 142134
rect 340826 102218 341062 102454
rect 341146 102218 341382 102454
rect 340826 101898 341062 102134
rect 341146 101898 341382 102134
rect 340826 62218 341062 62454
rect 341146 62218 341382 62454
rect 340826 61898 341062 62134
rect 341146 61898 341382 62134
rect 340826 22218 341062 22454
rect 341146 22218 341382 22454
rect 340826 21898 341062 22134
rect 341146 21898 341382 22134
rect 340826 -1542 341062 -1306
rect 341146 -1542 341382 -1306
rect 340826 -1862 341062 -1626
rect 341146 -1862 341382 -1626
rect 344546 665938 344782 666174
rect 344866 665938 345102 666174
rect 344546 665618 344782 665854
rect 344866 665618 345102 665854
rect 344546 625938 344782 626174
rect 344866 625938 345102 626174
rect 344546 625618 344782 625854
rect 344866 625618 345102 625854
rect 344546 585938 344782 586174
rect 344866 585938 345102 586174
rect 344546 585618 344782 585854
rect 344866 585618 345102 585854
rect 344546 545938 344782 546174
rect 344866 545938 345102 546174
rect 344546 545618 344782 545854
rect 344866 545618 345102 545854
rect 344546 505938 344782 506174
rect 344866 505938 345102 506174
rect 344546 505618 344782 505854
rect 344866 505618 345102 505854
rect 344546 465938 344782 466174
rect 344866 465938 345102 466174
rect 344546 465618 344782 465854
rect 344866 465618 345102 465854
rect 344546 425938 344782 426174
rect 344866 425938 345102 426174
rect 344546 425618 344782 425854
rect 344866 425618 345102 425854
rect 344546 385938 344782 386174
rect 344866 385938 345102 386174
rect 344546 385618 344782 385854
rect 344866 385618 345102 385854
rect 344546 345938 344782 346174
rect 344866 345938 345102 346174
rect 344546 345618 344782 345854
rect 344866 345618 345102 345854
rect 344546 305938 344782 306174
rect 344866 305938 345102 306174
rect 344546 305618 344782 305854
rect 344866 305618 345102 305854
rect 344546 265938 344782 266174
rect 344866 265938 345102 266174
rect 344546 265618 344782 265854
rect 344866 265618 345102 265854
rect 344546 225938 344782 226174
rect 344866 225938 345102 226174
rect 344546 225618 344782 225854
rect 344866 225618 345102 225854
rect 344546 185938 344782 186174
rect 344866 185938 345102 186174
rect 344546 185618 344782 185854
rect 344866 185618 345102 185854
rect 344546 145938 344782 146174
rect 344866 145938 345102 146174
rect 344546 145618 344782 145854
rect 344866 145618 345102 145854
rect 344546 105938 344782 106174
rect 344866 105938 345102 106174
rect 344546 105618 344782 105854
rect 344866 105618 345102 105854
rect 344546 65938 344782 66174
rect 344866 65938 345102 66174
rect 344546 65618 344782 65854
rect 344866 65618 345102 65854
rect 344546 25938 344782 26174
rect 344866 25938 345102 26174
rect 344546 25618 344782 25854
rect 344866 25618 345102 25854
rect 344546 -3462 344782 -3226
rect 344866 -3462 345102 -3226
rect 344546 -3782 344782 -3546
rect 344866 -3782 345102 -3546
rect 348266 669658 348502 669894
rect 348586 669658 348822 669894
rect 348266 669338 348502 669574
rect 348586 669338 348822 669574
rect 348266 629658 348502 629894
rect 348586 629658 348822 629894
rect 348266 629338 348502 629574
rect 348586 629338 348822 629574
rect 348266 589658 348502 589894
rect 348586 589658 348822 589894
rect 348266 589338 348502 589574
rect 348586 589338 348822 589574
rect 348266 549658 348502 549894
rect 348586 549658 348822 549894
rect 348266 549338 348502 549574
rect 348586 549338 348822 549574
rect 348266 509658 348502 509894
rect 348586 509658 348822 509894
rect 348266 509338 348502 509574
rect 348586 509338 348822 509574
rect 348266 469658 348502 469894
rect 348586 469658 348822 469894
rect 348266 469338 348502 469574
rect 348586 469338 348822 469574
rect 348266 429658 348502 429894
rect 348586 429658 348822 429894
rect 348266 429338 348502 429574
rect 348586 429338 348822 429574
rect 348266 389658 348502 389894
rect 348586 389658 348822 389894
rect 348266 389338 348502 389574
rect 348586 389338 348822 389574
rect 348266 349658 348502 349894
rect 348586 349658 348822 349894
rect 348266 349338 348502 349574
rect 348586 349338 348822 349574
rect 348266 309658 348502 309894
rect 348586 309658 348822 309894
rect 348266 309338 348502 309574
rect 348586 309338 348822 309574
rect 348266 269658 348502 269894
rect 348586 269658 348822 269894
rect 348266 269338 348502 269574
rect 348586 269338 348822 269574
rect 348266 229658 348502 229894
rect 348586 229658 348822 229894
rect 348266 229338 348502 229574
rect 348586 229338 348822 229574
rect 348266 189658 348502 189894
rect 348586 189658 348822 189894
rect 348266 189338 348502 189574
rect 348586 189338 348822 189574
rect 348266 149658 348502 149894
rect 348586 149658 348822 149894
rect 348266 149338 348502 149574
rect 348586 149338 348822 149574
rect 348266 109658 348502 109894
rect 348586 109658 348822 109894
rect 348266 109338 348502 109574
rect 348586 109338 348822 109574
rect 348266 69658 348502 69894
rect 348586 69658 348822 69894
rect 348266 69338 348502 69574
rect 348586 69338 348822 69574
rect 348266 29658 348502 29894
rect 348586 29658 348822 29894
rect 348266 29338 348502 29574
rect 348586 29338 348822 29574
rect 348266 -5382 348502 -5146
rect 348586 -5382 348822 -5146
rect 348266 -5702 348502 -5466
rect 348586 -5702 348822 -5466
rect 371986 710362 372222 710598
rect 372306 710362 372542 710598
rect 371986 710042 372222 710278
rect 372306 710042 372542 710278
rect 368266 708442 368502 708678
rect 368586 708442 368822 708678
rect 368266 708122 368502 708358
rect 368586 708122 368822 708358
rect 364546 706522 364782 706758
rect 364866 706522 365102 706758
rect 364546 706202 364782 706438
rect 364866 706202 365102 706438
rect 351986 673378 352222 673614
rect 352306 673378 352542 673614
rect 351986 673058 352222 673294
rect 352306 673058 352542 673294
rect 351986 633378 352222 633614
rect 352306 633378 352542 633614
rect 351986 633058 352222 633294
rect 352306 633058 352542 633294
rect 351986 593378 352222 593614
rect 352306 593378 352542 593614
rect 351986 593058 352222 593294
rect 352306 593058 352542 593294
rect 351986 553378 352222 553614
rect 352306 553378 352542 553614
rect 351986 553058 352222 553294
rect 352306 553058 352542 553294
rect 351986 513378 352222 513614
rect 352306 513378 352542 513614
rect 351986 513058 352222 513294
rect 352306 513058 352542 513294
rect 351986 473378 352222 473614
rect 352306 473378 352542 473614
rect 351986 473058 352222 473294
rect 352306 473058 352542 473294
rect 351986 433378 352222 433614
rect 352306 433378 352542 433614
rect 351986 433058 352222 433294
rect 352306 433058 352542 433294
rect 351986 393378 352222 393614
rect 352306 393378 352542 393614
rect 351986 393058 352222 393294
rect 352306 393058 352542 393294
rect 351986 353378 352222 353614
rect 352306 353378 352542 353614
rect 351986 353058 352222 353294
rect 352306 353058 352542 353294
rect 351986 313378 352222 313614
rect 352306 313378 352542 313614
rect 351986 313058 352222 313294
rect 352306 313058 352542 313294
rect 351986 273378 352222 273614
rect 352306 273378 352542 273614
rect 351986 273058 352222 273294
rect 352306 273058 352542 273294
rect 351986 233378 352222 233614
rect 352306 233378 352542 233614
rect 351986 233058 352222 233294
rect 352306 233058 352542 233294
rect 351986 193378 352222 193614
rect 352306 193378 352542 193614
rect 351986 193058 352222 193294
rect 352306 193058 352542 193294
rect 351986 153378 352222 153614
rect 352306 153378 352542 153614
rect 351986 153058 352222 153294
rect 352306 153058 352542 153294
rect 351986 113378 352222 113614
rect 352306 113378 352542 113614
rect 351986 113058 352222 113294
rect 352306 113058 352542 113294
rect 351986 73378 352222 73614
rect 352306 73378 352542 73614
rect 351986 73058 352222 73294
rect 352306 73058 352542 73294
rect 351986 33378 352222 33614
rect 352306 33378 352542 33614
rect 351986 33058 352222 33294
rect 352306 33058 352542 33294
rect 331986 -6342 332222 -6106
rect 332306 -6342 332542 -6106
rect 331986 -6662 332222 -6426
rect 332306 -6662 332542 -6426
rect 360826 704602 361062 704838
rect 361146 704602 361382 704838
rect 360826 704282 361062 704518
rect 361146 704282 361382 704518
rect 360826 682218 361062 682454
rect 361146 682218 361382 682454
rect 360826 681898 361062 682134
rect 361146 681898 361382 682134
rect 360826 642218 361062 642454
rect 361146 642218 361382 642454
rect 360826 641898 361062 642134
rect 361146 641898 361382 642134
rect 360826 602218 361062 602454
rect 361146 602218 361382 602454
rect 360826 601898 361062 602134
rect 361146 601898 361382 602134
rect 360826 562218 361062 562454
rect 361146 562218 361382 562454
rect 360826 561898 361062 562134
rect 361146 561898 361382 562134
rect 360826 522218 361062 522454
rect 361146 522218 361382 522454
rect 360826 521898 361062 522134
rect 361146 521898 361382 522134
rect 360826 482218 361062 482454
rect 361146 482218 361382 482454
rect 360826 481898 361062 482134
rect 361146 481898 361382 482134
rect 360826 442218 361062 442454
rect 361146 442218 361382 442454
rect 360826 441898 361062 442134
rect 361146 441898 361382 442134
rect 360826 402218 361062 402454
rect 361146 402218 361382 402454
rect 360826 401898 361062 402134
rect 361146 401898 361382 402134
rect 360826 362218 361062 362454
rect 361146 362218 361382 362454
rect 360826 361898 361062 362134
rect 361146 361898 361382 362134
rect 360826 322218 361062 322454
rect 361146 322218 361382 322454
rect 360826 321898 361062 322134
rect 361146 321898 361382 322134
rect 360826 282218 361062 282454
rect 361146 282218 361382 282454
rect 360826 281898 361062 282134
rect 361146 281898 361382 282134
rect 360826 242218 361062 242454
rect 361146 242218 361382 242454
rect 360826 241898 361062 242134
rect 361146 241898 361382 242134
rect 360826 202218 361062 202454
rect 361146 202218 361382 202454
rect 360826 201898 361062 202134
rect 361146 201898 361382 202134
rect 360826 162218 361062 162454
rect 361146 162218 361382 162454
rect 360826 161898 361062 162134
rect 361146 161898 361382 162134
rect 360826 122218 361062 122454
rect 361146 122218 361382 122454
rect 360826 121898 361062 122134
rect 361146 121898 361382 122134
rect 360826 82218 361062 82454
rect 361146 82218 361382 82454
rect 360826 81898 361062 82134
rect 361146 81898 361382 82134
rect 360826 42218 361062 42454
rect 361146 42218 361382 42454
rect 360826 41898 361062 42134
rect 361146 41898 361382 42134
rect 360826 2218 361062 2454
rect 361146 2218 361382 2454
rect 360826 1898 361062 2134
rect 361146 1898 361382 2134
rect 360826 -582 361062 -346
rect 361146 -582 361382 -346
rect 360826 -902 361062 -666
rect 361146 -902 361382 -666
rect 364546 685938 364782 686174
rect 364866 685938 365102 686174
rect 364546 685618 364782 685854
rect 364866 685618 365102 685854
rect 364546 645938 364782 646174
rect 364866 645938 365102 646174
rect 364546 645618 364782 645854
rect 364866 645618 365102 645854
rect 364546 605938 364782 606174
rect 364866 605938 365102 606174
rect 364546 605618 364782 605854
rect 364866 605618 365102 605854
rect 364546 565938 364782 566174
rect 364866 565938 365102 566174
rect 364546 565618 364782 565854
rect 364866 565618 365102 565854
rect 364546 525938 364782 526174
rect 364866 525938 365102 526174
rect 364546 525618 364782 525854
rect 364866 525618 365102 525854
rect 364546 485938 364782 486174
rect 364866 485938 365102 486174
rect 364546 485618 364782 485854
rect 364866 485618 365102 485854
rect 364546 445938 364782 446174
rect 364866 445938 365102 446174
rect 364546 445618 364782 445854
rect 364866 445618 365102 445854
rect 364546 405938 364782 406174
rect 364866 405938 365102 406174
rect 364546 405618 364782 405854
rect 364866 405618 365102 405854
rect 364546 365938 364782 366174
rect 364866 365938 365102 366174
rect 364546 365618 364782 365854
rect 364866 365618 365102 365854
rect 364546 325938 364782 326174
rect 364866 325938 365102 326174
rect 364546 325618 364782 325854
rect 364866 325618 365102 325854
rect 364546 285938 364782 286174
rect 364866 285938 365102 286174
rect 364546 285618 364782 285854
rect 364866 285618 365102 285854
rect 364546 245938 364782 246174
rect 364866 245938 365102 246174
rect 364546 245618 364782 245854
rect 364866 245618 365102 245854
rect 364546 205938 364782 206174
rect 364866 205938 365102 206174
rect 364546 205618 364782 205854
rect 364866 205618 365102 205854
rect 364546 165938 364782 166174
rect 364866 165938 365102 166174
rect 364546 165618 364782 165854
rect 364866 165618 365102 165854
rect 364546 125938 364782 126174
rect 364866 125938 365102 126174
rect 364546 125618 364782 125854
rect 364866 125618 365102 125854
rect 364546 85938 364782 86174
rect 364866 85938 365102 86174
rect 364546 85618 364782 85854
rect 364866 85618 365102 85854
rect 364546 45938 364782 46174
rect 364866 45938 365102 46174
rect 364546 45618 364782 45854
rect 364866 45618 365102 45854
rect 364546 5938 364782 6174
rect 364866 5938 365102 6174
rect 364546 5618 364782 5854
rect 364866 5618 365102 5854
rect 364546 -2502 364782 -2266
rect 364866 -2502 365102 -2266
rect 364546 -2822 364782 -2586
rect 364866 -2822 365102 -2586
rect 368266 689658 368502 689894
rect 368586 689658 368822 689894
rect 368266 689338 368502 689574
rect 368586 689338 368822 689574
rect 368266 649658 368502 649894
rect 368586 649658 368822 649894
rect 368266 649338 368502 649574
rect 368586 649338 368822 649574
rect 368266 609658 368502 609894
rect 368586 609658 368822 609894
rect 368266 609338 368502 609574
rect 368586 609338 368822 609574
rect 368266 569658 368502 569894
rect 368586 569658 368822 569894
rect 368266 569338 368502 569574
rect 368586 569338 368822 569574
rect 368266 529658 368502 529894
rect 368586 529658 368822 529894
rect 368266 529338 368502 529574
rect 368586 529338 368822 529574
rect 368266 489658 368502 489894
rect 368586 489658 368822 489894
rect 368266 489338 368502 489574
rect 368586 489338 368822 489574
rect 368266 449658 368502 449894
rect 368586 449658 368822 449894
rect 368266 449338 368502 449574
rect 368586 449338 368822 449574
rect 368266 409658 368502 409894
rect 368586 409658 368822 409894
rect 368266 409338 368502 409574
rect 368586 409338 368822 409574
rect 368266 369658 368502 369894
rect 368586 369658 368822 369894
rect 368266 369338 368502 369574
rect 368586 369338 368822 369574
rect 368266 329658 368502 329894
rect 368586 329658 368822 329894
rect 368266 329338 368502 329574
rect 368586 329338 368822 329574
rect 368266 289658 368502 289894
rect 368586 289658 368822 289894
rect 368266 289338 368502 289574
rect 368586 289338 368822 289574
rect 368266 249658 368502 249894
rect 368586 249658 368822 249894
rect 368266 249338 368502 249574
rect 368586 249338 368822 249574
rect 368266 209658 368502 209894
rect 368586 209658 368822 209894
rect 368266 209338 368502 209574
rect 368586 209338 368822 209574
rect 368266 169658 368502 169894
rect 368586 169658 368822 169894
rect 368266 169338 368502 169574
rect 368586 169338 368822 169574
rect 368266 129658 368502 129894
rect 368586 129658 368822 129894
rect 368266 129338 368502 129574
rect 368586 129338 368822 129574
rect 368266 89658 368502 89894
rect 368586 89658 368822 89894
rect 368266 89338 368502 89574
rect 368586 89338 368822 89574
rect 368266 49658 368502 49894
rect 368586 49658 368822 49894
rect 368266 49338 368502 49574
rect 368586 49338 368822 49574
rect 368266 9658 368502 9894
rect 368586 9658 368822 9894
rect 368266 9338 368502 9574
rect 368586 9338 368822 9574
rect 368266 -4422 368502 -4186
rect 368586 -4422 368822 -4186
rect 368266 -4742 368502 -4506
rect 368586 -4742 368822 -4506
rect 391986 711322 392222 711558
rect 392306 711322 392542 711558
rect 391986 711002 392222 711238
rect 392306 711002 392542 711238
rect 388266 709402 388502 709638
rect 388586 709402 388822 709638
rect 388266 709082 388502 709318
rect 388586 709082 388822 709318
rect 384546 707482 384782 707718
rect 384866 707482 385102 707718
rect 384546 707162 384782 707398
rect 384866 707162 385102 707398
rect 371986 693378 372222 693614
rect 372306 693378 372542 693614
rect 371986 693058 372222 693294
rect 372306 693058 372542 693294
rect 371986 653378 372222 653614
rect 372306 653378 372542 653614
rect 371986 653058 372222 653294
rect 372306 653058 372542 653294
rect 371986 613378 372222 613614
rect 372306 613378 372542 613614
rect 371986 613058 372222 613294
rect 372306 613058 372542 613294
rect 371986 573378 372222 573614
rect 372306 573378 372542 573614
rect 371986 573058 372222 573294
rect 372306 573058 372542 573294
rect 371986 533378 372222 533614
rect 372306 533378 372542 533614
rect 371986 533058 372222 533294
rect 372306 533058 372542 533294
rect 371986 493378 372222 493614
rect 372306 493378 372542 493614
rect 371986 493058 372222 493294
rect 372306 493058 372542 493294
rect 371986 453378 372222 453614
rect 372306 453378 372542 453614
rect 371986 453058 372222 453294
rect 372306 453058 372542 453294
rect 371986 413378 372222 413614
rect 372306 413378 372542 413614
rect 371986 413058 372222 413294
rect 372306 413058 372542 413294
rect 371986 373378 372222 373614
rect 372306 373378 372542 373614
rect 371986 373058 372222 373294
rect 372306 373058 372542 373294
rect 371986 333378 372222 333614
rect 372306 333378 372542 333614
rect 371986 333058 372222 333294
rect 372306 333058 372542 333294
rect 371986 293378 372222 293614
rect 372306 293378 372542 293614
rect 371986 293058 372222 293294
rect 372306 293058 372542 293294
rect 371986 253378 372222 253614
rect 372306 253378 372542 253614
rect 371986 253058 372222 253294
rect 372306 253058 372542 253294
rect 371986 213378 372222 213614
rect 372306 213378 372542 213614
rect 371986 213058 372222 213294
rect 372306 213058 372542 213294
rect 371986 173378 372222 173614
rect 372306 173378 372542 173614
rect 371986 173058 372222 173294
rect 372306 173058 372542 173294
rect 371986 133378 372222 133614
rect 372306 133378 372542 133614
rect 371986 133058 372222 133294
rect 372306 133058 372542 133294
rect 371986 93378 372222 93614
rect 372306 93378 372542 93614
rect 371986 93058 372222 93294
rect 372306 93058 372542 93294
rect 371986 53378 372222 53614
rect 372306 53378 372542 53614
rect 371986 53058 372222 53294
rect 372306 53058 372542 53294
rect 371986 13378 372222 13614
rect 372306 13378 372542 13614
rect 371986 13058 372222 13294
rect 372306 13058 372542 13294
rect 351986 -7302 352222 -7066
rect 352306 -7302 352542 -7066
rect 351986 -7622 352222 -7386
rect 352306 -7622 352542 -7386
rect 380826 705562 381062 705798
rect 381146 705562 381382 705798
rect 380826 705242 381062 705478
rect 381146 705242 381382 705478
rect 380826 662218 381062 662454
rect 381146 662218 381382 662454
rect 380826 661898 381062 662134
rect 381146 661898 381382 662134
rect 380826 622218 381062 622454
rect 381146 622218 381382 622454
rect 380826 621898 381062 622134
rect 381146 621898 381382 622134
rect 380826 582218 381062 582454
rect 381146 582218 381382 582454
rect 380826 581898 381062 582134
rect 381146 581898 381382 582134
rect 380826 542218 381062 542454
rect 381146 542218 381382 542454
rect 380826 541898 381062 542134
rect 381146 541898 381382 542134
rect 380826 502218 381062 502454
rect 381146 502218 381382 502454
rect 380826 501898 381062 502134
rect 381146 501898 381382 502134
rect 380826 462218 381062 462454
rect 381146 462218 381382 462454
rect 380826 461898 381062 462134
rect 381146 461898 381382 462134
rect 380826 422218 381062 422454
rect 381146 422218 381382 422454
rect 380826 421898 381062 422134
rect 381146 421898 381382 422134
rect 380826 382218 381062 382454
rect 381146 382218 381382 382454
rect 380826 381898 381062 382134
rect 381146 381898 381382 382134
rect 380826 342218 381062 342454
rect 381146 342218 381382 342454
rect 380826 341898 381062 342134
rect 381146 341898 381382 342134
rect 380826 302218 381062 302454
rect 381146 302218 381382 302454
rect 380826 301898 381062 302134
rect 381146 301898 381382 302134
rect 380826 262218 381062 262454
rect 381146 262218 381382 262454
rect 380826 261898 381062 262134
rect 381146 261898 381382 262134
rect 380826 222218 381062 222454
rect 381146 222218 381382 222454
rect 380826 221898 381062 222134
rect 381146 221898 381382 222134
rect 380826 182218 381062 182454
rect 381146 182218 381382 182454
rect 380826 181898 381062 182134
rect 381146 181898 381382 182134
rect 380826 142218 381062 142454
rect 381146 142218 381382 142454
rect 380826 141898 381062 142134
rect 381146 141898 381382 142134
rect 380826 102218 381062 102454
rect 381146 102218 381382 102454
rect 380826 101898 381062 102134
rect 381146 101898 381382 102134
rect 380826 62218 381062 62454
rect 381146 62218 381382 62454
rect 380826 61898 381062 62134
rect 381146 61898 381382 62134
rect 380826 22218 381062 22454
rect 381146 22218 381382 22454
rect 380826 21898 381062 22134
rect 381146 21898 381382 22134
rect 380826 -1542 381062 -1306
rect 381146 -1542 381382 -1306
rect 380826 -1862 381062 -1626
rect 381146 -1862 381382 -1626
rect 384546 665938 384782 666174
rect 384866 665938 385102 666174
rect 384546 665618 384782 665854
rect 384866 665618 385102 665854
rect 384546 625938 384782 626174
rect 384866 625938 385102 626174
rect 384546 625618 384782 625854
rect 384866 625618 385102 625854
rect 384546 585938 384782 586174
rect 384866 585938 385102 586174
rect 384546 585618 384782 585854
rect 384866 585618 385102 585854
rect 384546 545938 384782 546174
rect 384866 545938 385102 546174
rect 384546 545618 384782 545854
rect 384866 545618 385102 545854
rect 384546 505938 384782 506174
rect 384866 505938 385102 506174
rect 384546 505618 384782 505854
rect 384866 505618 385102 505854
rect 384546 465938 384782 466174
rect 384866 465938 385102 466174
rect 384546 465618 384782 465854
rect 384866 465618 385102 465854
rect 384546 425938 384782 426174
rect 384866 425938 385102 426174
rect 384546 425618 384782 425854
rect 384866 425618 385102 425854
rect 384546 385938 384782 386174
rect 384866 385938 385102 386174
rect 384546 385618 384782 385854
rect 384866 385618 385102 385854
rect 384546 345938 384782 346174
rect 384866 345938 385102 346174
rect 384546 345618 384782 345854
rect 384866 345618 385102 345854
rect 384546 305938 384782 306174
rect 384866 305938 385102 306174
rect 384546 305618 384782 305854
rect 384866 305618 385102 305854
rect 384546 265938 384782 266174
rect 384866 265938 385102 266174
rect 384546 265618 384782 265854
rect 384866 265618 385102 265854
rect 384546 225938 384782 226174
rect 384866 225938 385102 226174
rect 384546 225618 384782 225854
rect 384866 225618 385102 225854
rect 384546 185938 384782 186174
rect 384866 185938 385102 186174
rect 384546 185618 384782 185854
rect 384866 185618 385102 185854
rect 384546 145938 384782 146174
rect 384866 145938 385102 146174
rect 384546 145618 384782 145854
rect 384866 145618 385102 145854
rect 384546 105938 384782 106174
rect 384866 105938 385102 106174
rect 384546 105618 384782 105854
rect 384866 105618 385102 105854
rect 384546 65938 384782 66174
rect 384866 65938 385102 66174
rect 384546 65618 384782 65854
rect 384866 65618 385102 65854
rect 384546 25938 384782 26174
rect 384866 25938 385102 26174
rect 384546 25618 384782 25854
rect 384866 25618 385102 25854
rect 384546 -3462 384782 -3226
rect 384866 -3462 385102 -3226
rect 384546 -3782 384782 -3546
rect 384866 -3782 385102 -3546
rect 388266 669658 388502 669894
rect 388586 669658 388822 669894
rect 388266 669338 388502 669574
rect 388586 669338 388822 669574
rect 388266 629658 388502 629894
rect 388586 629658 388822 629894
rect 388266 629338 388502 629574
rect 388586 629338 388822 629574
rect 388266 589658 388502 589894
rect 388586 589658 388822 589894
rect 388266 589338 388502 589574
rect 388586 589338 388822 589574
rect 388266 549658 388502 549894
rect 388586 549658 388822 549894
rect 388266 549338 388502 549574
rect 388586 549338 388822 549574
rect 388266 509658 388502 509894
rect 388586 509658 388822 509894
rect 388266 509338 388502 509574
rect 388586 509338 388822 509574
rect 388266 469658 388502 469894
rect 388586 469658 388822 469894
rect 388266 469338 388502 469574
rect 388586 469338 388822 469574
rect 388266 429658 388502 429894
rect 388586 429658 388822 429894
rect 388266 429338 388502 429574
rect 388586 429338 388822 429574
rect 388266 389658 388502 389894
rect 388586 389658 388822 389894
rect 388266 389338 388502 389574
rect 388586 389338 388822 389574
rect 388266 349658 388502 349894
rect 388586 349658 388822 349894
rect 388266 349338 388502 349574
rect 388586 349338 388822 349574
rect 388266 309658 388502 309894
rect 388586 309658 388822 309894
rect 388266 309338 388502 309574
rect 388586 309338 388822 309574
rect 388266 269658 388502 269894
rect 388586 269658 388822 269894
rect 388266 269338 388502 269574
rect 388586 269338 388822 269574
rect 388266 229658 388502 229894
rect 388586 229658 388822 229894
rect 388266 229338 388502 229574
rect 388586 229338 388822 229574
rect 388266 189658 388502 189894
rect 388586 189658 388822 189894
rect 388266 189338 388502 189574
rect 388586 189338 388822 189574
rect 388266 149658 388502 149894
rect 388586 149658 388822 149894
rect 388266 149338 388502 149574
rect 388586 149338 388822 149574
rect 388266 109658 388502 109894
rect 388586 109658 388822 109894
rect 388266 109338 388502 109574
rect 388586 109338 388822 109574
rect 388266 69658 388502 69894
rect 388586 69658 388822 69894
rect 388266 69338 388502 69574
rect 388586 69338 388822 69574
rect 388266 29658 388502 29894
rect 388586 29658 388822 29894
rect 388266 29338 388502 29574
rect 388586 29338 388822 29574
rect 388266 -5382 388502 -5146
rect 388586 -5382 388822 -5146
rect 388266 -5702 388502 -5466
rect 388586 -5702 388822 -5466
rect 411986 710362 412222 710598
rect 412306 710362 412542 710598
rect 411986 710042 412222 710278
rect 412306 710042 412542 710278
rect 408266 708442 408502 708678
rect 408586 708442 408822 708678
rect 408266 708122 408502 708358
rect 408586 708122 408822 708358
rect 404546 706522 404782 706758
rect 404866 706522 405102 706758
rect 404546 706202 404782 706438
rect 404866 706202 405102 706438
rect 391986 673378 392222 673614
rect 392306 673378 392542 673614
rect 391986 673058 392222 673294
rect 392306 673058 392542 673294
rect 391986 633378 392222 633614
rect 392306 633378 392542 633614
rect 391986 633058 392222 633294
rect 392306 633058 392542 633294
rect 391986 593378 392222 593614
rect 392306 593378 392542 593614
rect 391986 593058 392222 593294
rect 392306 593058 392542 593294
rect 391986 553378 392222 553614
rect 392306 553378 392542 553614
rect 391986 553058 392222 553294
rect 392306 553058 392542 553294
rect 391986 513378 392222 513614
rect 392306 513378 392542 513614
rect 391986 513058 392222 513294
rect 392306 513058 392542 513294
rect 391986 473378 392222 473614
rect 392306 473378 392542 473614
rect 391986 473058 392222 473294
rect 392306 473058 392542 473294
rect 391986 433378 392222 433614
rect 392306 433378 392542 433614
rect 391986 433058 392222 433294
rect 392306 433058 392542 433294
rect 391986 393378 392222 393614
rect 392306 393378 392542 393614
rect 391986 393058 392222 393294
rect 392306 393058 392542 393294
rect 391986 353378 392222 353614
rect 392306 353378 392542 353614
rect 391986 353058 392222 353294
rect 392306 353058 392542 353294
rect 391986 313378 392222 313614
rect 392306 313378 392542 313614
rect 391986 313058 392222 313294
rect 392306 313058 392542 313294
rect 391986 273378 392222 273614
rect 392306 273378 392542 273614
rect 391986 273058 392222 273294
rect 392306 273058 392542 273294
rect 391986 233378 392222 233614
rect 392306 233378 392542 233614
rect 391986 233058 392222 233294
rect 392306 233058 392542 233294
rect 391986 193378 392222 193614
rect 392306 193378 392542 193614
rect 391986 193058 392222 193294
rect 392306 193058 392542 193294
rect 391986 153378 392222 153614
rect 392306 153378 392542 153614
rect 391986 153058 392222 153294
rect 392306 153058 392542 153294
rect 391986 113378 392222 113614
rect 392306 113378 392542 113614
rect 391986 113058 392222 113294
rect 392306 113058 392542 113294
rect 391986 73378 392222 73614
rect 392306 73378 392542 73614
rect 391986 73058 392222 73294
rect 392306 73058 392542 73294
rect 391986 33378 392222 33614
rect 392306 33378 392542 33614
rect 391986 33058 392222 33294
rect 392306 33058 392542 33294
rect 371986 -6342 372222 -6106
rect 372306 -6342 372542 -6106
rect 371986 -6662 372222 -6426
rect 372306 -6662 372542 -6426
rect 400826 704602 401062 704838
rect 401146 704602 401382 704838
rect 400826 704282 401062 704518
rect 401146 704282 401382 704518
rect 400826 682218 401062 682454
rect 401146 682218 401382 682454
rect 400826 681898 401062 682134
rect 401146 681898 401382 682134
rect 400826 642218 401062 642454
rect 401146 642218 401382 642454
rect 400826 641898 401062 642134
rect 401146 641898 401382 642134
rect 400826 602218 401062 602454
rect 401146 602218 401382 602454
rect 400826 601898 401062 602134
rect 401146 601898 401382 602134
rect 400826 562218 401062 562454
rect 401146 562218 401382 562454
rect 400826 561898 401062 562134
rect 401146 561898 401382 562134
rect 400826 522218 401062 522454
rect 401146 522218 401382 522454
rect 400826 521898 401062 522134
rect 401146 521898 401382 522134
rect 400826 482218 401062 482454
rect 401146 482218 401382 482454
rect 400826 481898 401062 482134
rect 401146 481898 401382 482134
rect 400826 442218 401062 442454
rect 401146 442218 401382 442454
rect 400826 441898 401062 442134
rect 401146 441898 401382 442134
rect 400826 402218 401062 402454
rect 401146 402218 401382 402454
rect 400826 401898 401062 402134
rect 401146 401898 401382 402134
rect 400826 362218 401062 362454
rect 401146 362218 401382 362454
rect 400826 361898 401062 362134
rect 401146 361898 401382 362134
rect 400826 322218 401062 322454
rect 401146 322218 401382 322454
rect 400826 321898 401062 322134
rect 401146 321898 401382 322134
rect 400826 282218 401062 282454
rect 401146 282218 401382 282454
rect 400826 281898 401062 282134
rect 401146 281898 401382 282134
rect 400826 242218 401062 242454
rect 401146 242218 401382 242454
rect 400826 241898 401062 242134
rect 401146 241898 401382 242134
rect 400826 202218 401062 202454
rect 401146 202218 401382 202454
rect 400826 201898 401062 202134
rect 401146 201898 401382 202134
rect 400826 162218 401062 162454
rect 401146 162218 401382 162454
rect 400826 161898 401062 162134
rect 401146 161898 401382 162134
rect 400826 122218 401062 122454
rect 401146 122218 401382 122454
rect 400826 121898 401062 122134
rect 401146 121898 401382 122134
rect 400826 82218 401062 82454
rect 401146 82218 401382 82454
rect 400826 81898 401062 82134
rect 401146 81898 401382 82134
rect 400826 42218 401062 42454
rect 401146 42218 401382 42454
rect 400826 41898 401062 42134
rect 401146 41898 401382 42134
rect 400826 2218 401062 2454
rect 401146 2218 401382 2454
rect 400826 1898 401062 2134
rect 401146 1898 401382 2134
rect 400826 -582 401062 -346
rect 401146 -582 401382 -346
rect 400826 -902 401062 -666
rect 401146 -902 401382 -666
rect 404546 685938 404782 686174
rect 404866 685938 405102 686174
rect 404546 685618 404782 685854
rect 404866 685618 405102 685854
rect 404546 645938 404782 646174
rect 404866 645938 405102 646174
rect 404546 645618 404782 645854
rect 404866 645618 405102 645854
rect 404546 605938 404782 606174
rect 404866 605938 405102 606174
rect 404546 605618 404782 605854
rect 404866 605618 405102 605854
rect 404546 565938 404782 566174
rect 404866 565938 405102 566174
rect 404546 565618 404782 565854
rect 404866 565618 405102 565854
rect 404546 525938 404782 526174
rect 404866 525938 405102 526174
rect 404546 525618 404782 525854
rect 404866 525618 405102 525854
rect 404546 485938 404782 486174
rect 404866 485938 405102 486174
rect 404546 485618 404782 485854
rect 404866 485618 405102 485854
rect 404546 445938 404782 446174
rect 404866 445938 405102 446174
rect 404546 445618 404782 445854
rect 404866 445618 405102 445854
rect 404546 405938 404782 406174
rect 404866 405938 405102 406174
rect 404546 405618 404782 405854
rect 404866 405618 405102 405854
rect 404546 365938 404782 366174
rect 404866 365938 405102 366174
rect 404546 365618 404782 365854
rect 404866 365618 405102 365854
rect 404546 325938 404782 326174
rect 404866 325938 405102 326174
rect 404546 325618 404782 325854
rect 404866 325618 405102 325854
rect 404546 285938 404782 286174
rect 404866 285938 405102 286174
rect 404546 285618 404782 285854
rect 404866 285618 405102 285854
rect 404546 245938 404782 246174
rect 404866 245938 405102 246174
rect 404546 245618 404782 245854
rect 404866 245618 405102 245854
rect 404546 205938 404782 206174
rect 404866 205938 405102 206174
rect 404546 205618 404782 205854
rect 404866 205618 405102 205854
rect 404546 165938 404782 166174
rect 404866 165938 405102 166174
rect 404546 165618 404782 165854
rect 404866 165618 405102 165854
rect 404546 125938 404782 126174
rect 404866 125938 405102 126174
rect 404546 125618 404782 125854
rect 404866 125618 405102 125854
rect 404546 85938 404782 86174
rect 404866 85938 405102 86174
rect 404546 85618 404782 85854
rect 404866 85618 405102 85854
rect 404546 45938 404782 46174
rect 404866 45938 405102 46174
rect 404546 45618 404782 45854
rect 404866 45618 405102 45854
rect 404546 5938 404782 6174
rect 404866 5938 405102 6174
rect 404546 5618 404782 5854
rect 404866 5618 405102 5854
rect 404546 -2502 404782 -2266
rect 404866 -2502 405102 -2266
rect 404546 -2822 404782 -2586
rect 404866 -2822 405102 -2586
rect 408266 689658 408502 689894
rect 408586 689658 408822 689894
rect 408266 689338 408502 689574
rect 408586 689338 408822 689574
rect 408266 649658 408502 649894
rect 408586 649658 408822 649894
rect 408266 649338 408502 649574
rect 408586 649338 408822 649574
rect 408266 609658 408502 609894
rect 408586 609658 408822 609894
rect 408266 609338 408502 609574
rect 408586 609338 408822 609574
rect 408266 569658 408502 569894
rect 408586 569658 408822 569894
rect 408266 569338 408502 569574
rect 408586 569338 408822 569574
rect 408266 529658 408502 529894
rect 408586 529658 408822 529894
rect 408266 529338 408502 529574
rect 408586 529338 408822 529574
rect 408266 489658 408502 489894
rect 408586 489658 408822 489894
rect 408266 489338 408502 489574
rect 408586 489338 408822 489574
rect 408266 449658 408502 449894
rect 408586 449658 408822 449894
rect 408266 449338 408502 449574
rect 408586 449338 408822 449574
rect 408266 409658 408502 409894
rect 408586 409658 408822 409894
rect 408266 409338 408502 409574
rect 408586 409338 408822 409574
rect 408266 369658 408502 369894
rect 408586 369658 408822 369894
rect 408266 369338 408502 369574
rect 408586 369338 408822 369574
rect 408266 329658 408502 329894
rect 408586 329658 408822 329894
rect 408266 329338 408502 329574
rect 408586 329338 408822 329574
rect 408266 289658 408502 289894
rect 408586 289658 408822 289894
rect 408266 289338 408502 289574
rect 408586 289338 408822 289574
rect 408266 249658 408502 249894
rect 408586 249658 408822 249894
rect 408266 249338 408502 249574
rect 408586 249338 408822 249574
rect 408266 209658 408502 209894
rect 408586 209658 408822 209894
rect 408266 209338 408502 209574
rect 408586 209338 408822 209574
rect 408266 169658 408502 169894
rect 408586 169658 408822 169894
rect 408266 169338 408502 169574
rect 408586 169338 408822 169574
rect 408266 129658 408502 129894
rect 408586 129658 408822 129894
rect 408266 129338 408502 129574
rect 408586 129338 408822 129574
rect 408266 89658 408502 89894
rect 408586 89658 408822 89894
rect 408266 89338 408502 89574
rect 408586 89338 408822 89574
rect 408266 49658 408502 49894
rect 408586 49658 408822 49894
rect 408266 49338 408502 49574
rect 408586 49338 408822 49574
rect 408266 9658 408502 9894
rect 408586 9658 408822 9894
rect 408266 9338 408502 9574
rect 408586 9338 408822 9574
rect 408266 -4422 408502 -4186
rect 408586 -4422 408822 -4186
rect 408266 -4742 408502 -4506
rect 408586 -4742 408822 -4506
rect 431986 711322 432222 711558
rect 432306 711322 432542 711558
rect 431986 711002 432222 711238
rect 432306 711002 432542 711238
rect 428266 709402 428502 709638
rect 428586 709402 428822 709638
rect 428266 709082 428502 709318
rect 428586 709082 428822 709318
rect 424546 707482 424782 707718
rect 424866 707482 425102 707718
rect 424546 707162 424782 707398
rect 424866 707162 425102 707398
rect 411986 693378 412222 693614
rect 412306 693378 412542 693614
rect 411986 693058 412222 693294
rect 412306 693058 412542 693294
rect 411986 653378 412222 653614
rect 412306 653378 412542 653614
rect 411986 653058 412222 653294
rect 412306 653058 412542 653294
rect 411986 613378 412222 613614
rect 412306 613378 412542 613614
rect 411986 613058 412222 613294
rect 412306 613058 412542 613294
rect 411986 573378 412222 573614
rect 412306 573378 412542 573614
rect 411986 573058 412222 573294
rect 412306 573058 412542 573294
rect 411986 533378 412222 533614
rect 412306 533378 412542 533614
rect 411986 533058 412222 533294
rect 412306 533058 412542 533294
rect 411986 493378 412222 493614
rect 412306 493378 412542 493614
rect 411986 493058 412222 493294
rect 412306 493058 412542 493294
rect 411986 453378 412222 453614
rect 412306 453378 412542 453614
rect 411986 453058 412222 453294
rect 412306 453058 412542 453294
rect 411986 413378 412222 413614
rect 412306 413378 412542 413614
rect 411986 413058 412222 413294
rect 412306 413058 412542 413294
rect 411986 373378 412222 373614
rect 412306 373378 412542 373614
rect 411986 373058 412222 373294
rect 412306 373058 412542 373294
rect 411986 333378 412222 333614
rect 412306 333378 412542 333614
rect 411986 333058 412222 333294
rect 412306 333058 412542 333294
rect 411986 293378 412222 293614
rect 412306 293378 412542 293614
rect 411986 293058 412222 293294
rect 412306 293058 412542 293294
rect 411986 253378 412222 253614
rect 412306 253378 412542 253614
rect 411986 253058 412222 253294
rect 412306 253058 412542 253294
rect 411986 213378 412222 213614
rect 412306 213378 412542 213614
rect 411986 213058 412222 213294
rect 412306 213058 412542 213294
rect 411986 173378 412222 173614
rect 412306 173378 412542 173614
rect 411986 173058 412222 173294
rect 412306 173058 412542 173294
rect 411986 133378 412222 133614
rect 412306 133378 412542 133614
rect 411986 133058 412222 133294
rect 412306 133058 412542 133294
rect 411986 93378 412222 93614
rect 412306 93378 412542 93614
rect 411986 93058 412222 93294
rect 412306 93058 412542 93294
rect 411986 53378 412222 53614
rect 412306 53378 412542 53614
rect 411986 53058 412222 53294
rect 412306 53058 412542 53294
rect 411986 13378 412222 13614
rect 412306 13378 412542 13614
rect 411986 13058 412222 13294
rect 412306 13058 412542 13294
rect 391986 -7302 392222 -7066
rect 392306 -7302 392542 -7066
rect 391986 -7622 392222 -7386
rect 392306 -7622 392542 -7386
rect 420826 705562 421062 705798
rect 421146 705562 421382 705798
rect 420826 705242 421062 705478
rect 421146 705242 421382 705478
rect 420826 662218 421062 662454
rect 421146 662218 421382 662454
rect 420826 661898 421062 662134
rect 421146 661898 421382 662134
rect 420826 622218 421062 622454
rect 421146 622218 421382 622454
rect 420826 621898 421062 622134
rect 421146 621898 421382 622134
rect 420826 582218 421062 582454
rect 421146 582218 421382 582454
rect 420826 581898 421062 582134
rect 421146 581898 421382 582134
rect 420826 542218 421062 542454
rect 421146 542218 421382 542454
rect 420826 541898 421062 542134
rect 421146 541898 421382 542134
rect 420826 502218 421062 502454
rect 421146 502218 421382 502454
rect 420826 501898 421062 502134
rect 421146 501898 421382 502134
rect 420826 462218 421062 462454
rect 421146 462218 421382 462454
rect 420826 461898 421062 462134
rect 421146 461898 421382 462134
rect 420826 422218 421062 422454
rect 421146 422218 421382 422454
rect 420826 421898 421062 422134
rect 421146 421898 421382 422134
rect 420826 382218 421062 382454
rect 421146 382218 421382 382454
rect 420826 381898 421062 382134
rect 421146 381898 421382 382134
rect 420826 342218 421062 342454
rect 421146 342218 421382 342454
rect 420826 341898 421062 342134
rect 421146 341898 421382 342134
rect 420826 302218 421062 302454
rect 421146 302218 421382 302454
rect 420826 301898 421062 302134
rect 421146 301898 421382 302134
rect 420826 262218 421062 262454
rect 421146 262218 421382 262454
rect 420826 261898 421062 262134
rect 421146 261898 421382 262134
rect 420826 222218 421062 222454
rect 421146 222218 421382 222454
rect 420826 221898 421062 222134
rect 421146 221898 421382 222134
rect 420826 182218 421062 182454
rect 421146 182218 421382 182454
rect 420826 181898 421062 182134
rect 421146 181898 421382 182134
rect 420826 142218 421062 142454
rect 421146 142218 421382 142454
rect 420826 141898 421062 142134
rect 421146 141898 421382 142134
rect 420826 102218 421062 102454
rect 421146 102218 421382 102454
rect 420826 101898 421062 102134
rect 421146 101898 421382 102134
rect 420826 62218 421062 62454
rect 421146 62218 421382 62454
rect 420826 61898 421062 62134
rect 421146 61898 421382 62134
rect 420826 22218 421062 22454
rect 421146 22218 421382 22454
rect 420826 21898 421062 22134
rect 421146 21898 421382 22134
rect 420826 -1542 421062 -1306
rect 421146 -1542 421382 -1306
rect 420826 -1862 421062 -1626
rect 421146 -1862 421382 -1626
rect 424546 665938 424782 666174
rect 424866 665938 425102 666174
rect 424546 665618 424782 665854
rect 424866 665618 425102 665854
rect 424546 625938 424782 626174
rect 424866 625938 425102 626174
rect 424546 625618 424782 625854
rect 424866 625618 425102 625854
rect 424546 585938 424782 586174
rect 424866 585938 425102 586174
rect 424546 585618 424782 585854
rect 424866 585618 425102 585854
rect 424546 545938 424782 546174
rect 424866 545938 425102 546174
rect 424546 545618 424782 545854
rect 424866 545618 425102 545854
rect 424546 505938 424782 506174
rect 424866 505938 425102 506174
rect 424546 505618 424782 505854
rect 424866 505618 425102 505854
rect 424546 465938 424782 466174
rect 424866 465938 425102 466174
rect 424546 465618 424782 465854
rect 424866 465618 425102 465854
rect 424546 425938 424782 426174
rect 424866 425938 425102 426174
rect 424546 425618 424782 425854
rect 424866 425618 425102 425854
rect 424546 385938 424782 386174
rect 424866 385938 425102 386174
rect 424546 385618 424782 385854
rect 424866 385618 425102 385854
rect 424546 345938 424782 346174
rect 424866 345938 425102 346174
rect 424546 345618 424782 345854
rect 424866 345618 425102 345854
rect 424546 305938 424782 306174
rect 424866 305938 425102 306174
rect 424546 305618 424782 305854
rect 424866 305618 425102 305854
rect 424546 265938 424782 266174
rect 424866 265938 425102 266174
rect 424546 265618 424782 265854
rect 424866 265618 425102 265854
rect 424546 225938 424782 226174
rect 424866 225938 425102 226174
rect 424546 225618 424782 225854
rect 424866 225618 425102 225854
rect 424546 185938 424782 186174
rect 424866 185938 425102 186174
rect 424546 185618 424782 185854
rect 424866 185618 425102 185854
rect 424546 145938 424782 146174
rect 424866 145938 425102 146174
rect 424546 145618 424782 145854
rect 424866 145618 425102 145854
rect 424546 105938 424782 106174
rect 424866 105938 425102 106174
rect 424546 105618 424782 105854
rect 424866 105618 425102 105854
rect 424546 65938 424782 66174
rect 424866 65938 425102 66174
rect 424546 65618 424782 65854
rect 424866 65618 425102 65854
rect 424546 25938 424782 26174
rect 424866 25938 425102 26174
rect 424546 25618 424782 25854
rect 424866 25618 425102 25854
rect 424546 -3462 424782 -3226
rect 424866 -3462 425102 -3226
rect 424546 -3782 424782 -3546
rect 424866 -3782 425102 -3546
rect 428266 669658 428502 669894
rect 428586 669658 428822 669894
rect 428266 669338 428502 669574
rect 428586 669338 428822 669574
rect 428266 629658 428502 629894
rect 428586 629658 428822 629894
rect 428266 629338 428502 629574
rect 428586 629338 428822 629574
rect 428266 589658 428502 589894
rect 428586 589658 428822 589894
rect 428266 589338 428502 589574
rect 428586 589338 428822 589574
rect 428266 549658 428502 549894
rect 428586 549658 428822 549894
rect 428266 549338 428502 549574
rect 428586 549338 428822 549574
rect 428266 509658 428502 509894
rect 428586 509658 428822 509894
rect 428266 509338 428502 509574
rect 428586 509338 428822 509574
rect 428266 469658 428502 469894
rect 428586 469658 428822 469894
rect 428266 469338 428502 469574
rect 428586 469338 428822 469574
rect 428266 429658 428502 429894
rect 428586 429658 428822 429894
rect 428266 429338 428502 429574
rect 428586 429338 428822 429574
rect 428266 389658 428502 389894
rect 428586 389658 428822 389894
rect 428266 389338 428502 389574
rect 428586 389338 428822 389574
rect 428266 349658 428502 349894
rect 428586 349658 428822 349894
rect 428266 349338 428502 349574
rect 428586 349338 428822 349574
rect 428266 309658 428502 309894
rect 428586 309658 428822 309894
rect 428266 309338 428502 309574
rect 428586 309338 428822 309574
rect 428266 269658 428502 269894
rect 428586 269658 428822 269894
rect 428266 269338 428502 269574
rect 428586 269338 428822 269574
rect 428266 229658 428502 229894
rect 428586 229658 428822 229894
rect 428266 229338 428502 229574
rect 428586 229338 428822 229574
rect 428266 189658 428502 189894
rect 428586 189658 428822 189894
rect 428266 189338 428502 189574
rect 428586 189338 428822 189574
rect 428266 149658 428502 149894
rect 428586 149658 428822 149894
rect 428266 149338 428502 149574
rect 428586 149338 428822 149574
rect 428266 109658 428502 109894
rect 428586 109658 428822 109894
rect 428266 109338 428502 109574
rect 428586 109338 428822 109574
rect 428266 69658 428502 69894
rect 428586 69658 428822 69894
rect 428266 69338 428502 69574
rect 428586 69338 428822 69574
rect 428266 29658 428502 29894
rect 428586 29658 428822 29894
rect 428266 29338 428502 29574
rect 428586 29338 428822 29574
rect 428266 -5382 428502 -5146
rect 428586 -5382 428822 -5146
rect 428266 -5702 428502 -5466
rect 428586 -5702 428822 -5466
rect 451986 710362 452222 710598
rect 452306 710362 452542 710598
rect 451986 710042 452222 710278
rect 452306 710042 452542 710278
rect 448266 708442 448502 708678
rect 448586 708442 448822 708678
rect 448266 708122 448502 708358
rect 448586 708122 448822 708358
rect 444546 706522 444782 706758
rect 444866 706522 445102 706758
rect 444546 706202 444782 706438
rect 444866 706202 445102 706438
rect 431986 673378 432222 673614
rect 432306 673378 432542 673614
rect 431986 673058 432222 673294
rect 432306 673058 432542 673294
rect 431986 633378 432222 633614
rect 432306 633378 432542 633614
rect 431986 633058 432222 633294
rect 432306 633058 432542 633294
rect 431986 593378 432222 593614
rect 432306 593378 432542 593614
rect 431986 593058 432222 593294
rect 432306 593058 432542 593294
rect 431986 553378 432222 553614
rect 432306 553378 432542 553614
rect 431986 553058 432222 553294
rect 432306 553058 432542 553294
rect 431986 513378 432222 513614
rect 432306 513378 432542 513614
rect 431986 513058 432222 513294
rect 432306 513058 432542 513294
rect 431986 473378 432222 473614
rect 432306 473378 432542 473614
rect 431986 473058 432222 473294
rect 432306 473058 432542 473294
rect 431986 433378 432222 433614
rect 432306 433378 432542 433614
rect 431986 433058 432222 433294
rect 432306 433058 432542 433294
rect 431986 393378 432222 393614
rect 432306 393378 432542 393614
rect 431986 393058 432222 393294
rect 432306 393058 432542 393294
rect 431986 353378 432222 353614
rect 432306 353378 432542 353614
rect 431986 353058 432222 353294
rect 432306 353058 432542 353294
rect 431986 313378 432222 313614
rect 432306 313378 432542 313614
rect 431986 313058 432222 313294
rect 432306 313058 432542 313294
rect 431986 273378 432222 273614
rect 432306 273378 432542 273614
rect 431986 273058 432222 273294
rect 432306 273058 432542 273294
rect 431986 233378 432222 233614
rect 432306 233378 432542 233614
rect 431986 233058 432222 233294
rect 432306 233058 432542 233294
rect 431986 193378 432222 193614
rect 432306 193378 432542 193614
rect 431986 193058 432222 193294
rect 432306 193058 432542 193294
rect 431986 153378 432222 153614
rect 432306 153378 432542 153614
rect 431986 153058 432222 153294
rect 432306 153058 432542 153294
rect 431986 113378 432222 113614
rect 432306 113378 432542 113614
rect 431986 113058 432222 113294
rect 432306 113058 432542 113294
rect 431986 73378 432222 73614
rect 432306 73378 432542 73614
rect 431986 73058 432222 73294
rect 432306 73058 432542 73294
rect 431986 33378 432222 33614
rect 432306 33378 432542 33614
rect 431986 33058 432222 33294
rect 432306 33058 432542 33294
rect 411986 -6342 412222 -6106
rect 412306 -6342 412542 -6106
rect 411986 -6662 412222 -6426
rect 412306 -6662 412542 -6426
rect 440826 704602 441062 704838
rect 441146 704602 441382 704838
rect 440826 704282 441062 704518
rect 441146 704282 441382 704518
rect 440826 682218 441062 682454
rect 441146 682218 441382 682454
rect 440826 681898 441062 682134
rect 441146 681898 441382 682134
rect 440826 642218 441062 642454
rect 441146 642218 441382 642454
rect 440826 641898 441062 642134
rect 441146 641898 441382 642134
rect 440826 602218 441062 602454
rect 441146 602218 441382 602454
rect 440826 601898 441062 602134
rect 441146 601898 441382 602134
rect 440826 562218 441062 562454
rect 441146 562218 441382 562454
rect 440826 561898 441062 562134
rect 441146 561898 441382 562134
rect 440826 522218 441062 522454
rect 441146 522218 441382 522454
rect 440826 521898 441062 522134
rect 441146 521898 441382 522134
rect 440826 482218 441062 482454
rect 441146 482218 441382 482454
rect 440826 481898 441062 482134
rect 441146 481898 441382 482134
rect 440826 442218 441062 442454
rect 441146 442218 441382 442454
rect 440826 441898 441062 442134
rect 441146 441898 441382 442134
rect 440826 402218 441062 402454
rect 441146 402218 441382 402454
rect 440826 401898 441062 402134
rect 441146 401898 441382 402134
rect 440826 362218 441062 362454
rect 441146 362218 441382 362454
rect 440826 361898 441062 362134
rect 441146 361898 441382 362134
rect 440826 322218 441062 322454
rect 441146 322218 441382 322454
rect 440826 321898 441062 322134
rect 441146 321898 441382 322134
rect 440826 282218 441062 282454
rect 441146 282218 441382 282454
rect 440826 281898 441062 282134
rect 441146 281898 441382 282134
rect 440826 242218 441062 242454
rect 441146 242218 441382 242454
rect 440826 241898 441062 242134
rect 441146 241898 441382 242134
rect 440826 202218 441062 202454
rect 441146 202218 441382 202454
rect 440826 201898 441062 202134
rect 441146 201898 441382 202134
rect 440826 162218 441062 162454
rect 441146 162218 441382 162454
rect 440826 161898 441062 162134
rect 441146 161898 441382 162134
rect 440826 122218 441062 122454
rect 441146 122218 441382 122454
rect 440826 121898 441062 122134
rect 441146 121898 441382 122134
rect 440826 82218 441062 82454
rect 441146 82218 441382 82454
rect 440826 81898 441062 82134
rect 441146 81898 441382 82134
rect 440826 42218 441062 42454
rect 441146 42218 441382 42454
rect 440826 41898 441062 42134
rect 441146 41898 441382 42134
rect 440826 2218 441062 2454
rect 441146 2218 441382 2454
rect 440826 1898 441062 2134
rect 441146 1898 441382 2134
rect 440826 -582 441062 -346
rect 441146 -582 441382 -346
rect 440826 -902 441062 -666
rect 441146 -902 441382 -666
rect 444546 685938 444782 686174
rect 444866 685938 445102 686174
rect 444546 685618 444782 685854
rect 444866 685618 445102 685854
rect 444546 645938 444782 646174
rect 444866 645938 445102 646174
rect 444546 645618 444782 645854
rect 444866 645618 445102 645854
rect 444546 605938 444782 606174
rect 444866 605938 445102 606174
rect 444546 605618 444782 605854
rect 444866 605618 445102 605854
rect 444546 565938 444782 566174
rect 444866 565938 445102 566174
rect 444546 565618 444782 565854
rect 444866 565618 445102 565854
rect 444546 525938 444782 526174
rect 444866 525938 445102 526174
rect 444546 525618 444782 525854
rect 444866 525618 445102 525854
rect 444546 485938 444782 486174
rect 444866 485938 445102 486174
rect 444546 485618 444782 485854
rect 444866 485618 445102 485854
rect 444546 445938 444782 446174
rect 444866 445938 445102 446174
rect 444546 445618 444782 445854
rect 444866 445618 445102 445854
rect 444546 405938 444782 406174
rect 444866 405938 445102 406174
rect 444546 405618 444782 405854
rect 444866 405618 445102 405854
rect 444546 365938 444782 366174
rect 444866 365938 445102 366174
rect 444546 365618 444782 365854
rect 444866 365618 445102 365854
rect 444546 325938 444782 326174
rect 444866 325938 445102 326174
rect 444546 325618 444782 325854
rect 444866 325618 445102 325854
rect 444546 285938 444782 286174
rect 444866 285938 445102 286174
rect 444546 285618 444782 285854
rect 444866 285618 445102 285854
rect 444546 245938 444782 246174
rect 444866 245938 445102 246174
rect 444546 245618 444782 245854
rect 444866 245618 445102 245854
rect 444546 205938 444782 206174
rect 444866 205938 445102 206174
rect 444546 205618 444782 205854
rect 444866 205618 445102 205854
rect 444546 165938 444782 166174
rect 444866 165938 445102 166174
rect 444546 165618 444782 165854
rect 444866 165618 445102 165854
rect 444546 125938 444782 126174
rect 444866 125938 445102 126174
rect 444546 125618 444782 125854
rect 444866 125618 445102 125854
rect 444546 85938 444782 86174
rect 444866 85938 445102 86174
rect 444546 85618 444782 85854
rect 444866 85618 445102 85854
rect 444546 45938 444782 46174
rect 444866 45938 445102 46174
rect 444546 45618 444782 45854
rect 444866 45618 445102 45854
rect 444546 5938 444782 6174
rect 444866 5938 445102 6174
rect 444546 5618 444782 5854
rect 444866 5618 445102 5854
rect 444546 -2502 444782 -2266
rect 444866 -2502 445102 -2266
rect 444546 -2822 444782 -2586
rect 444866 -2822 445102 -2586
rect 448266 689658 448502 689894
rect 448586 689658 448822 689894
rect 448266 689338 448502 689574
rect 448586 689338 448822 689574
rect 448266 649658 448502 649894
rect 448586 649658 448822 649894
rect 448266 649338 448502 649574
rect 448586 649338 448822 649574
rect 448266 609658 448502 609894
rect 448586 609658 448822 609894
rect 448266 609338 448502 609574
rect 448586 609338 448822 609574
rect 448266 569658 448502 569894
rect 448586 569658 448822 569894
rect 448266 569338 448502 569574
rect 448586 569338 448822 569574
rect 448266 529658 448502 529894
rect 448586 529658 448822 529894
rect 448266 529338 448502 529574
rect 448586 529338 448822 529574
rect 448266 489658 448502 489894
rect 448586 489658 448822 489894
rect 448266 489338 448502 489574
rect 448586 489338 448822 489574
rect 448266 449658 448502 449894
rect 448586 449658 448822 449894
rect 448266 449338 448502 449574
rect 448586 449338 448822 449574
rect 448266 409658 448502 409894
rect 448586 409658 448822 409894
rect 448266 409338 448502 409574
rect 448586 409338 448822 409574
rect 448266 369658 448502 369894
rect 448586 369658 448822 369894
rect 448266 369338 448502 369574
rect 448586 369338 448822 369574
rect 448266 329658 448502 329894
rect 448586 329658 448822 329894
rect 448266 329338 448502 329574
rect 448586 329338 448822 329574
rect 448266 289658 448502 289894
rect 448586 289658 448822 289894
rect 448266 289338 448502 289574
rect 448586 289338 448822 289574
rect 448266 249658 448502 249894
rect 448586 249658 448822 249894
rect 448266 249338 448502 249574
rect 448586 249338 448822 249574
rect 448266 209658 448502 209894
rect 448586 209658 448822 209894
rect 448266 209338 448502 209574
rect 448586 209338 448822 209574
rect 448266 169658 448502 169894
rect 448586 169658 448822 169894
rect 448266 169338 448502 169574
rect 448586 169338 448822 169574
rect 448266 129658 448502 129894
rect 448586 129658 448822 129894
rect 448266 129338 448502 129574
rect 448586 129338 448822 129574
rect 448266 89658 448502 89894
rect 448586 89658 448822 89894
rect 448266 89338 448502 89574
rect 448586 89338 448822 89574
rect 448266 49658 448502 49894
rect 448586 49658 448822 49894
rect 448266 49338 448502 49574
rect 448586 49338 448822 49574
rect 448266 9658 448502 9894
rect 448586 9658 448822 9894
rect 448266 9338 448502 9574
rect 448586 9338 448822 9574
rect 448266 -4422 448502 -4186
rect 448586 -4422 448822 -4186
rect 448266 -4742 448502 -4506
rect 448586 -4742 448822 -4506
rect 471986 711322 472222 711558
rect 472306 711322 472542 711558
rect 471986 711002 472222 711238
rect 472306 711002 472542 711238
rect 468266 709402 468502 709638
rect 468586 709402 468822 709638
rect 468266 709082 468502 709318
rect 468586 709082 468822 709318
rect 464546 707482 464782 707718
rect 464866 707482 465102 707718
rect 464546 707162 464782 707398
rect 464866 707162 465102 707398
rect 451986 693378 452222 693614
rect 452306 693378 452542 693614
rect 451986 693058 452222 693294
rect 452306 693058 452542 693294
rect 451986 653378 452222 653614
rect 452306 653378 452542 653614
rect 451986 653058 452222 653294
rect 452306 653058 452542 653294
rect 451986 613378 452222 613614
rect 452306 613378 452542 613614
rect 451986 613058 452222 613294
rect 452306 613058 452542 613294
rect 451986 573378 452222 573614
rect 452306 573378 452542 573614
rect 451986 573058 452222 573294
rect 452306 573058 452542 573294
rect 451986 533378 452222 533614
rect 452306 533378 452542 533614
rect 451986 533058 452222 533294
rect 452306 533058 452542 533294
rect 451986 493378 452222 493614
rect 452306 493378 452542 493614
rect 451986 493058 452222 493294
rect 452306 493058 452542 493294
rect 451986 453378 452222 453614
rect 452306 453378 452542 453614
rect 451986 453058 452222 453294
rect 452306 453058 452542 453294
rect 451986 413378 452222 413614
rect 452306 413378 452542 413614
rect 451986 413058 452222 413294
rect 452306 413058 452542 413294
rect 451986 373378 452222 373614
rect 452306 373378 452542 373614
rect 451986 373058 452222 373294
rect 452306 373058 452542 373294
rect 451986 333378 452222 333614
rect 452306 333378 452542 333614
rect 451986 333058 452222 333294
rect 452306 333058 452542 333294
rect 451986 293378 452222 293614
rect 452306 293378 452542 293614
rect 451986 293058 452222 293294
rect 452306 293058 452542 293294
rect 451986 253378 452222 253614
rect 452306 253378 452542 253614
rect 451986 253058 452222 253294
rect 452306 253058 452542 253294
rect 451986 213378 452222 213614
rect 452306 213378 452542 213614
rect 451986 213058 452222 213294
rect 452306 213058 452542 213294
rect 451986 173378 452222 173614
rect 452306 173378 452542 173614
rect 451986 173058 452222 173294
rect 452306 173058 452542 173294
rect 451986 133378 452222 133614
rect 452306 133378 452542 133614
rect 451986 133058 452222 133294
rect 452306 133058 452542 133294
rect 451986 93378 452222 93614
rect 452306 93378 452542 93614
rect 451986 93058 452222 93294
rect 452306 93058 452542 93294
rect 451986 53378 452222 53614
rect 452306 53378 452542 53614
rect 451986 53058 452222 53294
rect 452306 53058 452542 53294
rect 451986 13378 452222 13614
rect 452306 13378 452542 13614
rect 451986 13058 452222 13294
rect 452306 13058 452542 13294
rect 431986 -7302 432222 -7066
rect 432306 -7302 432542 -7066
rect 431986 -7622 432222 -7386
rect 432306 -7622 432542 -7386
rect 460826 705562 461062 705798
rect 461146 705562 461382 705798
rect 460826 705242 461062 705478
rect 461146 705242 461382 705478
rect 460826 662218 461062 662454
rect 461146 662218 461382 662454
rect 460826 661898 461062 662134
rect 461146 661898 461382 662134
rect 460826 622218 461062 622454
rect 461146 622218 461382 622454
rect 460826 621898 461062 622134
rect 461146 621898 461382 622134
rect 460826 582218 461062 582454
rect 461146 582218 461382 582454
rect 460826 581898 461062 582134
rect 461146 581898 461382 582134
rect 460826 542218 461062 542454
rect 461146 542218 461382 542454
rect 460826 541898 461062 542134
rect 461146 541898 461382 542134
rect 460826 502218 461062 502454
rect 461146 502218 461382 502454
rect 460826 501898 461062 502134
rect 461146 501898 461382 502134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 422218 461062 422454
rect 461146 422218 461382 422454
rect 460826 421898 461062 422134
rect 461146 421898 461382 422134
rect 460826 382218 461062 382454
rect 461146 382218 461382 382454
rect 460826 381898 461062 382134
rect 461146 381898 461382 382134
rect 460826 342218 461062 342454
rect 461146 342218 461382 342454
rect 460826 341898 461062 342134
rect 461146 341898 461382 342134
rect 460826 302218 461062 302454
rect 461146 302218 461382 302454
rect 460826 301898 461062 302134
rect 461146 301898 461382 302134
rect 460826 262218 461062 262454
rect 461146 262218 461382 262454
rect 460826 261898 461062 262134
rect 461146 261898 461382 262134
rect 460826 222218 461062 222454
rect 461146 222218 461382 222454
rect 460826 221898 461062 222134
rect 461146 221898 461382 222134
rect 460826 182218 461062 182454
rect 461146 182218 461382 182454
rect 460826 181898 461062 182134
rect 461146 181898 461382 182134
rect 460826 142218 461062 142454
rect 461146 142218 461382 142454
rect 460826 141898 461062 142134
rect 461146 141898 461382 142134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 62218 461062 62454
rect 461146 62218 461382 62454
rect 460826 61898 461062 62134
rect 461146 61898 461382 62134
rect 460826 22218 461062 22454
rect 461146 22218 461382 22454
rect 460826 21898 461062 22134
rect 461146 21898 461382 22134
rect 460826 -1542 461062 -1306
rect 461146 -1542 461382 -1306
rect 460826 -1862 461062 -1626
rect 461146 -1862 461382 -1626
rect 464546 665938 464782 666174
rect 464866 665938 465102 666174
rect 464546 665618 464782 665854
rect 464866 665618 465102 665854
rect 464546 625938 464782 626174
rect 464866 625938 465102 626174
rect 464546 625618 464782 625854
rect 464866 625618 465102 625854
rect 464546 585938 464782 586174
rect 464866 585938 465102 586174
rect 464546 585618 464782 585854
rect 464866 585618 465102 585854
rect 464546 545938 464782 546174
rect 464866 545938 465102 546174
rect 464546 545618 464782 545854
rect 464866 545618 465102 545854
rect 464546 505938 464782 506174
rect 464866 505938 465102 506174
rect 464546 505618 464782 505854
rect 464866 505618 465102 505854
rect 464546 465938 464782 466174
rect 464866 465938 465102 466174
rect 464546 465618 464782 465854
rect 464866 465618 465102 465854
rect 464546 425938 464782 426174
rect 464866 425938 465102 426174
rect 464546 425618 464782 425854
rect 464866 425618 465102 425854
rect 464546 385938 464782 386174
rect 464866 385938 465102 386174
rect 464546 385618 464782 385854
rect 464866 385618 465102 385854
rect 464546 345938 464782 346174
rect 464866 345938 465102 346174
rect 464546 345618 464782 345854
rect 464866 345618 465102 345854
rect 464546 305938 464782 306174
rect 464866 305938 465102 306174
rect 464546 305618 464782 305854
rect 464866 305618 465102 305854
rect 464546 265938 464782 266174
rect 464866 265938 465102 266174
rect 464546 265618 464782 265854
rect 464866 265618 465102 265854
rect 464546 225938 464782 226174
rect 464866 225938 465102 226174
rect 464546 225618 464782 225854
rect 464866 225618 465102 225854
rect 464546 185938 464782 186174
rect 464866 185938 465102 186174
rect 464546 185618 464782 185854
rect 464866 185618 465102 185854
rect 464546 145938 464782 146174
rect 464866 145938 465102 146174
rect 464546 145618 464782 145854
rect 464866 145618 465102 145854
rect 464546 105938 464782 106174
rect 464866 105938 465102 106174
rect 464546 105618 464782 105854
rect 464866 105618 465102 105854
rect 464546 65938 464782 66174
rect 464866 65938 465102 66174
rect 464546 65618 464782 65854
rect 464866 65618 465102 65854
rect 464546 25938 464782 26174
rect 464866 25938 465102 26174
rect 464546 25618 464782 25854
rect 464866 25618 465102 25854
rect 464546 -3462 464782 -3226
rect 464866 -3462 465102 -3226
rect 464546 -3782 464782 -3546
rect 464866 -3782 465102 -3546
rect 468266 669658 468502 669894
rect 468586 669658 468822 669894
rect 468266 669338 468502 669574
rect 468586 669338 468822 669574
rect 468266 629658 468502 629894
rect 468586 629658 468822 629894
rect 468266 629338 468502 629574
rect 468586 629338 468822 629574
rect 468266 589658 468502 589894
rect 468586 589658 468822 589894
rect 468266 589338 468502 589574
rect 468586 589338 468822 589574
rect 468266 549658 468502 549894
rect 468586 549658 468822 549894
rect 468266 549338 468502 549574
rect 468586 549338 468822 549574
rect 468266 509658 468502 509894
rect 468586 509658 468822 509894
rect 468266 509338 468502 509574
rect 468586 509338 468822 509574
rect 468266 469658 468502 469894
rect 468586 469658 468822 469894
rect 468266 469338 468502 469574
rect 468586 469338 468822 469574
rect 468266 429658 468502 429894
rect 468586 429658 468822 429894
rect 468266 429338 468502 429574
rect 468586 429338 468822 429574
rect 468266 389658 468502 389894
rect 468586 389658 468822 389894
rect 468266 389338 468502 389574
rect 468586 389338 468822 389574
rect 468266 349658 468502 349894
rect 468586 349658 468822 349894
rect 468266 349338 468502 349574
rect 468586 349338 468822 349574
rect 468266 309658 468502 309894
rect 468586 309658 468822 309894
rect 468266 309338 468502 309574
rect 468586 309338 468822 309574
rect 468266 269658 468502 269894
rect 468586 269658 468822 269894
rect 468266 269338 468502 269574
rect 468586 269338 468822 269574
rect 468266 229658 468502 229894
rect 468586 229658 468822 229894
rect 468266 229338 468502 229574
rect 468586 229338 468822 229574
rect 468266 189658 468502 189894
rect 468586 189658 468822 189894
rect 468266 189338 468502 189574
rect 468586 189338 468822 189574
rect 468266 149658 468502 149894
rect 468586 149658 468822 149894
rect 468266 149338 468502 149574
rect 468586 149338 468822 149574
rect 468266 109658 468502 109894
rect 468586 109658 468822 109894
rect 468266 109338 468502 109574
rect 468586 109338 468822 109574
rect 468266 69658 468502 69894
rect 468586 69658 468822 69894
rect 468266 69338 468502 69574
rect 468586 69338 468822 69574
rect 468266 29658 468502 29894
rect 468586 29658 468822 29894
rect 468266 29338 468502 29574
rect 468586 29338 468822 29574
rect 468266 -5382 468502 -5146
rect 468586 -5382 468822 -5146
rect 468266 -5702 468502 -5466
rect 468586 -5702 468822 -5466
rect 491986 710362 492222 710598
rect 492306 710362 492542 710598
rect 491986 710042 492222 710278
rect 492306 710042 492542 710278
rect 488266 708442 488502 708678
rect 488586 708442 488822 708678
rect 488266 708122 488502 708358
rect 488586 708122 488822 708358
rect 484546 706522 484782 706758
rect 484866 706522 485102 706758
rect 484546 706202 484782 706438
rect 484866 706202 485102 706438
rect 471986 673378 472222 673614
rect 472306 673378 472542 673614
rect 471986 673058 472222 673294
rect 472306 673058 472542 673294
rect 471986 633378 472222 633614
rect 472306 633378 472542 633614
rect 471986 633058 472222 633294
rect 472306 633058 472542 633294
rect 471986 593378 472222 593614
rect 472306 593378 472542 593614
rect 471986 593058 472222 593294
rect 472306 593058 472542 593294
rect 471986 553378 472222 553614
rect 472306 553378 472542 553614
rect 471986 553058 472222 553294
rect 472306 553058 472542 553294
rect 471986 513378 472222 513614
rect 472306 513378 472542 513614
rect 471986 513058 472222 513294
rect 472306 513058 472542 513294
rect 471986 473378 472222 473614
rect 472306 473378 472542 473614
rect 471986 473058 472222 473294
rect 472306 473058 472542 473294
rect 471986 433378 472222 433614
rect 472306 433378 472542 433614
rect 471986 433058 472222 433294
rect 472306 433058 472542 433294
rect 471986 393378 472222 393614
rect 472306 393378 472542 393614
rect 471986 393058 472222 393294
rect 472306 393058 472542 393294
rect 471986 353378 472222 353614
rect 472306 353378 472542 353614
rect 471986 353058 472222 353294
rect 472306 353058 472542 353294
rect 471986 313378 472222 313614
rect 472306 313378 472542 313614
rect 471986 313058 472222 313294
rect 472306 313058 472542 313294
rect 471986 273378 472222 273614
rect 472306 273378 472542 273614
rect 471986 273058 472222 273294
rect 472306 273058 472542 273294
rect 471986 233378 472222 233614
rect 472306 233378 472542 233614
rect 471986 233058 472222 233294
rect 472306 233058 472542 233294
rect 471986 193378 472222 193614
rect 472306 193378 472542 193614
rect 471986 193058 472222 193294
rect 472306 193058 472542 193294
rect 471986 153378 472222 153614
rect 472306 153378 472542 153614
rect 471986 153058 472222 153294
rect 472306 153058 472542 153294
rect 471986 113378 472222 113614
rect 472306 113378 472542 113614
rect 471986 113058 472222 113294
rect 472306 113058 472542 113294
rect 471986 73378 472222 73614
rect 472306 73378 472542 73614
rect 471986 73058 472222 73294
rect 472306 73058 472542 73294
rect 471986 33378 472222 33614
rect 472306 33378 472542 33614
rect 471986 33058 472222 33294
rect 472306 33058 472542 33294
rect 451986 -6342 452222 -6106
rect 452306 -6342 452542 -6106
rect 451986 -6662 452222 -6426
rect 452306 -6662 452542 -6426
rect 480826 704602 481062 704838
rect 481146 704602 481382 704838
rect 480826 704282 481062 704518
rect 481146 704282 481382 704518
rect 480826 682218 481062 682454
rect 481146 682218 481382 682454
rect 480826 681898 481062 682134
rect 481146 681898 481382 682134
rect 480826 642218 481062 642454
rect 481146 642218 481382 642454
rect 480826 641898 481062 642134
rect 481146 641898 481382 642134
rect 480826 602218 481062 602454
rect 481146 602218 481382 602454
rect 480826 601898 481062 602134
rect 481146 601898 481382 602134
rect 480826 562218 481062 562454
rect 481146 562218 481382 562454
rect 480826 561898 481062 562134
rect 481146 561898 481382 562134
rect 480826 522218 481062 522454
rect 481146 522218 481382 522454
rect 480826 521898 481062 522134
rect 481146 521898 481382 522134
rect 480826 482218 481062 482454
rect 481146 482218 481382 482454
rect 480826 481898 481062 482134
rect 481146 481898 481382 482134
rect 480826 442218 481062 442454
rect 481146 442218 481382 442454
rect 480826 441898 481062 442134
rect 481146 441898 481382 442134
rect 480826 402218 481062 402454
rect 481146 402218 481382 402454
rect 480826 401898 481062 402134
rect 481146 401898 481382 402134
rect 480826 362218 481062 362454
rect 481146 362218 481382 362454
rect 480826 361898 481062 362134
rect 481146 361898 481382 362134
rect 480826 322218 481062 322454
rect 481146 322218 481382 322454
rect 480826 321898 481062 322134
rect 481146 321898 481382 322134
rect 480826 282218 481062 282454
rect 481146 282218 481382 282454
rect 480826 281898 481062 282134
rect 481146 281898 481382 282134
rect 480826 242218 481062 242454
rect 481146 242218 481382 242454
rect 480826 241898 481062 242134
rect 481146 241898 481382 242134
rect 480826 202218 481062 202454
rect 481146 202218 481382 202454
rect 480826 201898 481062 202134
rect 481146 201898 481382 202134
rect 480826 162218 481062 162454
rect 481146 162218 481382 162454
rect 480826 161898 481062 162134
rect 481146 161898 481382 162134
rect 480826 122218 481062 122454
rect 481146 122218 481382 122454
rect 480826 121898 481062 122134
rect 481146 121898 481382 122134
rect 480826 82218 481062 82454
rect 481146 82218 481382 82454
rect 480826 81898 481062 82134
rect 481146 81898 481382 82134
rect 480826 42218 481062 42454
rect 481146 42218 481382 42454
rect 480826 41898 481062 42134
rect 481146 41898 481382 42134
rect 480826 2218 481062 2454
rect 481146 2218 481382 2454
rect 480826 1898 481062 2134
rect 481146 1898 481382 2134
rect 480826 -582 481062 -346
rect 481146 -582 481382 -346
rect 480826 -902 481062 -666
rect 481146 -902 481382 -666
rect 484546 685938 484782 686174
rect 484866 685938 485102 686174
rect 484546 685618 484782 685854
rect 484866 685618 485102 685854
rect 484546 645938 484782 646174
rect 484866 645938 485102 646174
rect 484546 645618 484782 645854
rect 484866 645618 485102 645854
rect 484546 605938 484782 606174
rect 484866 605938 485102 606174
rect 484546 605618 484782 605854
rect 484866 605618 485102 605854
rect 484546 565938 484782 566174
rect 484866 565938 485102 566174
rect 484546 565618 484782 565854
rect 484866 565618 485102 565854
rect 484546 525938 484782 526174
rect 484866 525938 485102 526174
rect 484546 525618 484782 525854
rect 484866 525618 485102 525854
rect 484546 485938 484782 486174
rect 484866 485938 485102 486174
rect 484546 485618 484782 485854
rect 484866 485618 485102 485854
rect 484546 445938 484782 446174
rect 484866 445938 485102 446174
rect 484546 445618 484782 445854
rect 484866 445618 485102 445854
rect 484546 405938 484782 406174
rect 484866 405938 485102 406174
rect 484546 405618 484782 405854
rect 484866 405618 485102 405854
rect 484546 365938 484782 366174
rect 484866 365938 485102 366174
rect 484546 365618 484782 365854
rect 484866 365618 485102 365854
rect 484546 325938 484782 326174
rect 484866 325938 485102 326174
rect 484546 325618 484782 325854
rect 484866 325618 485102 325854
rect 484546 285938 484782 286174
rect 484866 285938 485102 286174
rect 484546 285618 484782 285854
rect 484866 285618 485102 285854
rect 484546 245938 484782 246174
rect 484866 245938 485102 246174
rect 484546 245618 484782 245854
rect 484866 245618 485102 245854
rect 484546 205938 484782 206174
rect 484866 205938 485102 206174
rect 484546 205618 484782 205854
rect 484866 205618 485102 205854
rect 484546 165938 484782 166174
rect 484866 165938 485102 166174
rect 484546 165618 484782 165854
rect 484866 165618 485102 165854
rect 484546 125938 484782 126174
rect 484866 125938 485102 126174
rect 484546 125618 484782 125854
rect 484866 125618 485102 125854
rect 484546 85938 484782 86174
rect 484866 85938 485102 86174
rect 484546 85618 484782 85854
rect 484866 85618 485102 85854
rect 484546 45938 484782 46174
rect 484866 45938 485102 46174
rect 484546 45618 484782 45854
rect 484866 45618 485102 45854
rect 484546 5938 484782 6174
rect 484866 5938 485102 6174
rect 484546 5618 484782 5854
rect 484866 5618 485102 5854
rect 484546 -2502 484782 -2266
rect 484866 -2502 485102 -2266
rect 484546 -2822 484782 -2586
rect 484866 -2822 485102 -2586
rect 488266 689658 488502 689894
rect 488586 689658 488822 689894
rect 488266 689338 488502 689574
rect 488586 689338 488822 689574
rect 488266 649658 488502 649894
rect 488586 649658 488822 649894
rect 488266 649338 488502 649574
rect 488586 649338 488822 649574
rect 488266 609658 488502 609894
rect 488586 609658 488822 609894
rect 488266 609338 488502 609574
rect 488586 609338 488822 609574
rect 488266 569658 488502 569894
rect 488586 569658 488822 569894
rect 488266 569338 488502 569574
rect 488586 569338 488822 569574
rect 488266 529658 488502 529894
rect 488586 529658 488822 529894
rect 488266 529338 488502 529574
rect 488586 529338 488822 529574
rect 488266 489658 488502 489894
rect 488586 489658 488822 489894
rect 488266 489338 488502 489574
rect 488586 489338 488822 489574
rect 488266 449658 488502 449894
rect 488586 449658 488822 449894
rect 488266 449338 488502 449574
rect 488586 449338 488822 449574
rect 488266 409658 488502 409894
rect 488586 409658 488822 409894
rect 488266 409338 488502 409574
rect 488586 409338 488822 409574
rect 488266 369658 488502 369894
rect 488586 369658 488822 369894
rect 488266 369338 488502 369574
rect 488586 369338 488822 369574
rect 488266 329658 488502 329894
rect 488586 329658 488822 329894
rect 488266 329338 488502 329574
rect 488586 329338 488822 329574
rect 488266 289658 488502 289894
rect 488586 289658 488822 289894
rect 488266 289338 488502 289574
rect 488586 289338 488822 289574
rect 488266 249658 488502 249894
rect 488586 249658 488822 249894
rect 488266 249338 488502 249574
rect 488586 249338 488822 249574
rect 488266 209658 488502 209894
rect 488586 209658 488822 209894
rect 488266 209338 488502 209574
rect 488586 209338 488822 209574
rect 488266 169658 488502 169894
rect 488586 169658 488822 169894
rect 488266 169338 488502 169574
rect 488586 169338 488822 169574
rect 488266 129658 488502 129894
rect 488586 129658 488822 129894
rect 488266 129338 488502 129574
rect 488586 129338 488822 129574
rect 488266 89658 488502 89894
rect 488586 89658 488822 89894
rect 488266 89338 488502 89574
rect 488586 89338 488822 89574
rect 488266 49658 488502 49894
rect 488586 49658 488822 49894
rect 488266 49338 488502 49574
rect 488586 49338 488822 49574
rect 488266 9658 488502 9894
rect 488586 9658 488822 9894
rect 488266 9338 488502 9574
rect 488586 9338 488822 9574
rect 488266 -4422 488502 -4186
rect 488586 -4422 488822 -4186
rect 488266 -4742 488502 -4506
rect 488586 -4742 488822 -4506
rect 511986 711322 512222 711558
rect 512306 711322 512542 711558
rect 511986 711002 512222 711238
rect 512306 711002 512542 711238
rect 508266 709402 508502 709638
rect 508586 709402 508822 709638
rect 508266 709082 508502 709318
rect 508586 709082 508822 709318
rect 504546 707482 504782 707718
rect 504866 707482 505102 707718
rect 504546 707162 504782 707398
rect 504866 707162 505102 707398
rect 491986 693378 492222 693614
rect 492306 693378 492542 693614
rect 491986 693058 492222 693294
rect 492306 693058 492542 693294
rect 491986 653378 492222 653614
rect 492306 653378 492542 653614
rect 491986 653058 492222 653294
rect 492306 653058 492542 653294
rect 491986 613378 492222 613614
rect 492306 613378 492542 613614
rect 491986 613058 492222 613294
rect 492306 613058 492542 613294
rect 491986 573378 492222 573614
rect 492306 573378 492542 573614
rect 491986 573058 492222 573294
rect 492306 573058 492542 573294
rect 491986 533378 492222 533614
rect 492306 533378 492542 533614
rect 491986 533058 492222 533294
rect 492306 533058 492542 533294
rect 491986 493378 492222 493614
rect 492306 493378 492542 493614
rect 491986 493058 492222 493294
rect 492306 493058 492542 493294
rect 491986 453378 492222 453614
rect 492306 453378 492542 453614
rect 491986 453058 492222 453294
rect 492306 453058 492542 453294
rect 491986 413378 492222 413614
rect 492306 413378 492542 413614
rect 491986 413058 492222 413294
rect 492306 413058 492542 413294
rect 491986 373378 492222 373614
rect 492306 373378 492542 373614
rect 491986 373058 492222 373294
rect 492306 373058 492542 373294
rect 491986 333378 492222 333614
rect 492306 333378 492542 333614
rect 491986 333058 492222 333294
rect 492306 333058 492542 333294
rect 491986 293378 492222 293614
rect 492306 293378 492542 293614
rect 491986 293058 492222 293294
rect 492306 293058 492542 293294
rect 491986 253378 492222 253614
rect 492306 253378 492542 253614
rect 491986 253058 492222 253294
rect 492306 253058 492542 253294
rect 491986 213378 492222 213614
rect 492306 213378 492542 213614
rect 491986 213058 492222 213294
rect 492306 213058 492542 213294
rect 491986 173378 492222 173614
rect 492306 173378 492542 173614
rect 491986 173058 492222 173294
rect 492306 173058 492542 173294
rect 491986 133378 492222 133614
rect 492306 133378 492542 133614
rect 491986 133058 492222 133294
rect 492306 133058 492542 133294
rect 491986 93378 492222 93614
rect 492306 93378 492542 93614
rect 491986 93058 492222 93294
rect 492306 93058 492542 93294
rect 491986 53378 492222 53614
rect 492306 53378 492542 53614
rect 491986 53058 492222 53294
rect 492306 53058 492542 53294
rect 491986 13378 492222 13614
rect 492306 13378 492542 13614
rect 491986 13058 492222 13294
rect 492306 13058 492542 13294
rect 471986 -7302 472222 -7066
rect 472306 -7302 472542 -7066
rect 471986 -7622 472222 -7386
rect 472306 -7622 472542 -7386
rect 500826 705562 501062 705798
rect 501146 705562 501382 705798
rect 500826 705242 501062 705478
rect 501146 705242 501382 705478
rect 500826 662218 501062 662454
rect 501146 662218 501382 662454
rect 500826 661898 501062 662134
rect 501146 661898 501382 662134
rect 500826 622218 501062 622454
rect 501146 622218 501382 622454
rect 500826 621898 501062 622134
rect 501146 621898 501382 622134
rect 500826 582218 501062 582454
rect 501146 582218 501382 582454
rect 500826 581898 501062 582134
rect 501146 581898 501382 582134
rect 500826 542218 501062 542454
rect 501146 542218 501382 542454
rect 500826 541898 501062 542134
rect 501146 541898 501382 542134
rect 500826 502218 501062 502454
rect 501146 502218 501382 502454
rect 500826 501898 501062 502134
rect 501146 501898 501382 502134
rect 500826 462218 501062 462454
rect 501146 462218 501382 462454
rect 500826 461898 501062 462134
rect 501146 461898 501382 462134
rect 500826 422218 501062 422454
rect 501146 422218 501382 422454
rect 500826 421898 501062 422134
rect 501146 421898 501382 422134
rect 500826 382218 501062 382454
rect 501146 382218 501382 382454
rect 500826 381898 501062 382134
rect 501146 381898 501382 382134
rect 500826 342218 501062 342454
rect 501146 342218 501382 342454
rect 500826 341898 501062 342134
rect 501146 341898 501382 342134
rect 500826 302218 501062 302454
rect 501146 302218 501382 302454
rect 500826 301898 501062 302134
rect 501146 301898 501382 302134
rect 500826 262218 501062 262454
rect 501146 262218 501382 262454
rect 500826 261898 501062 262134
rect 501146 261898 501382 262134
rect 500826 222218 501062 222454
rect 501146 222218 501382 222454
rect 500826 221898 501062 222134
rect 501146 221898 501382 222134
rect 500826 182218 501062 182454
rect 501146 182218 501382 182454
rect 500826 181898 501062 182134
rect 501146 181898 501382 182134
rect 500826 142218 501062 142454
rect 501146 142218 501382 142454
rect 500826 141898 501062 142134
rect 501146 141898 501382 142134
rect 500826 102218 501062 102454
rect 501146 102218 501382 102454
rect 500826 101898 501062 102134
rect 501146 101898 501382 102134
rect 500826 62218 501062 62454
rect 501146 62218 501382 62454
rect 500826 61898 501062 62134
rect 501146 61898 501382 62134
rect 500826 22218 501062 22454
rect 501146 22218 501382 22454
rect 500826 21898 501062 22134
rect 501146 21898 501382 22134
rect 500826 -1542 501062 -1306
rect 501146 -1542 501382 -1306
rect 500826 -1862 501062 -1626
rect 501146 -1862 501382 -1626
rect 504546 665938 504782 666174
rect 504866 665938 505102 666174
rect 504546 665618 504782 665854
rect 504866 665618 505102 665854
rect 504546 625938 504782 626174
rect 504866 625938 505102 626174
rect 504546 625618 504782 625854
rect 504866 625618 505102 625854
rect 504546 585938 504782 586174
rect 504866 585938 505102 586174
rect 504546 585618 504782 585854
rect 504866 585618 505102 585854
rect 504546 545938 504782 546174
rect 504866 545938 505102 546174
rect 504546 545618 504782 545854
rect 504866 545618 505102 545854
rect 504546 505938 504782 506174
rect 504866 505938 505102 506174
rect 504546 505618 504782 505854
rect 504866 505618 505102 505854
rect 504546 465938 504782 466174
rect 504866 465938 505102 466174
rect 504546 465618 504782 465854
rect 504866 465618 505102 465854
rect 504546 425938 504782 426174
rect 504866 425938 505102 426174
rect 504546 425618 504782 425854
rect 504866 425618 505102 425854
rect 504546 385938 504782 386174
rect 504866 385938 505102 386174
rect 504546 385618 504782 385854
rect 504866 385618 505102 385854
rect 504546 345938 504782 346174
rect 504866 345938 505102 346174
rect 504546 345618 504782 345854
rect 504866 345618 505102 345854
rect 504546 305938 504782 306174
rect 504866 305938 505102 306174
rect 504546 305618 504782 305854
rect 504866 305618 505102 305854
rect 504546 265938 504782 266174
rect 504866 265938 505102 266174
rect 504546 265618 504782 265854
rect 504866 265618 505102 265854
rect 504546 225938 504782 226174
rect 504866 225938 505102 226174
rect 504546 225618 504782 225854
rect 504866 225618 505102 225854
rect 504546 185938 504782 186174
rect 504866 185938 505102 186174
rect 504546 185618 504782 185854
rect 504866 185618 505102 185854
rect 504546 145938 504782 146174
rect 504866 145938 505102 146174
rect 504546 145618 504782 145854
rect 504866 145618 505102 145854
rect 504546 105938 504782 106174
rect 504866 105938 505102 106174
rect 504546 105618 504782 105854
rect 504866 105618 505102 105854
rect 504546 65938 504782 66174
rect 504866 65938 505102 66174
rect 504546 65618 504782 65854
rect 504866 65618 505102 65854
rect 504546 25938 504782 26174
rect 504866 25938 505102 26174
rect 504546 25618 504782 25854
rect 504866 25618 505102 25854
rect 504546 -3462 504782 -3226
rect 504866 -3462 505102 -3226
rect 504546 -3782 504782 -3546
rect 504866 -3782 505102 -3546
rect 508266 669658 508502 669894
rect 508586 669658 508822 669894
rect 508266 669338 508502 669574
rect 508586 669338 508822 669574
rect 508266 629658 508502 629894
rect 508586 629658 508822 629894
rect 508266 629338 508502 629574
rect 508586 629338 508822 629574
rect 508266 589658 508502 589894
rect 508586 589658 508822 589894
rect 508266 589338 508502 589574
rect 508586 589338 508822 589574
rect 508266 549658 508502 549894
rect 508586 549658 508822 549894
rect 508266 549338 508502 549574
rect 508586 549338 508822 549574
rect 508266 509658 508502 509894
rect 508586 509658 508822 509894
rect 508266 509338 508502 509574
rect 508586 509338 508822 509574
rect 508266 469658 508502 469894
rect 508586 469658 508822 469894
rect 508266 469338 508502 469574
rect 508586 469338 508822 469574
rect 508266 429658 508502 429894
rect 508586 429658 508822 429894
rect 508266 429338 508502 429574
rect 508586 429338 508822 429574
rect 508266 389658 508502 389894
rect 508586 389658 508822 389894
rect 508266 389338 508502 389574
rect 508586 389338 508822 389574
rect 508266 349658 508502 349894
rect 508586 349658 508822 349894
rect 508266 349338 508502 349574
rect 508586 349338 508822 349574
rect 508266 309658 508502 309894
rect 508586 309658 508822 309894
rect 508266 309338 508502 309574
rect 508586 309338 508822 309574
rect 508266 269658 508502 269894
rect 508586 269658 508822 269894
rect 508266 269338 508502 269574
rect 508586 269338 508822 269574
rect 508266 229658 508502 229894
rect 508586 229658 508822 229894
rect 508266 229338 508502 229574
rect 508586 229338 508822 229574
rect 508266 189658 508502 189894
rect 508586 189658 508822 189894
rect 508266 189338 508502 189574
rect 508586 189338 508822 189574
rect 508266 149658 508502 149894
rect 508586 149658 508822 149894
rect 508266 149338 508502 149574
rect 508586 149338 508822 149574
rect 508266 109658 508502 109894
rect 508586 109658 508822 109894
rect 508266 109338 508502 109574
rect 508586 109338 508822 109574
rect 508266 69658 508502 69894
rect 508586 69658 508822 69894
rect 508266 69338 508502 69574
rect 508586 69338 508822 69574
rect 508266 29658 508502 29894
rect 508586 29658 508822 29894
rect 508266 29338 508502 29574
rect 508586 29338 508822 29574
rect 508266 -5382 508502 -5146
rect 508586 -5382 508822 -5146
rect 508266 -5702 508502 -5466
rect 508586 -5702 508822 -5466
rect 531986 710362 532222 710598
rect 532306 710362 532542 710598
rect 531986 710042 532222 710278
rect 532306 710042 532542 710278
rect 528266 708442 528502 708678
rect 528586 708442 528822 708678
rect 528266 708122 528502 708358
rect 528586 708122 528822 708358
rect 524546 706522 524782 706758
rect 524866 706522 525102 706758
rect 524546 706202 524782 706438
rect 524866 706202 525102 706438
rect 511986 673378 512222 673614
rect 512306 673378 512542 673614
rect 511986 673058 512222 673294
rect 512306 673058 512542 673294
rect 511986 633378 512222 633614
rect 512306 633378 512542 633614
rect 511986 633058 512222 633294
rect 512306 633058 512542 633294
rect 511986 593378 512222 593614
rect 512306 593378 512542 593614
rect 511986 593058 512222 593294
rect 512306 593058 512542 593294
rect 511986 553378 512222 553614
rect 512306 553378 512542 553614
rect 511986 553058 512222 553294
rect 512306 553058 512542 553294
rect 511986 513378 512222 513614
rect 512306 513378 512542 513614
rect 511986 513058 512222 513294
rect 512306 513058 512542 513294
rect 511986 473378 512222 473614
rect 512306 473378 512542 473614
rect 511986 473058 512222 473294
rect 512306 473058 512542 473294
rect 511986 433378 512222 433614
rect 512306 433378 512542 433614
rect 511986 433058 512222 433294
rect 512306 433058 512542 433294
rect 511986 393378 512222 393614
rect 512306 393378 512542 393614
rect 511986 393058 512222 393294
rect 512306 393058 512542 393294
rect 511986 353378 512222 353614
rect 512306 353378 512542 353614
rect 511986 353058 512222 353294
rect 512306 353058 512542 353294
rect 511986 313378 512222 313614
rect 512306 313378 512542 313614
rect 511986 313058 512222 313294
rect 512306 313058 512542 313294
rect 511986 273378 512222 273614
rect 512306 273378 512542 273614
rect 511986 273058 512222 273294
rect 512306 273058 512542 273294
rect 511986 233378 512222 233614
rect 512306 233378 512542 233614
rect 511986 233058 512222 233294
rect 512306 233058 512542 233294
rect 511986 193378 512222 193614
rect 512306 193378 512542 193614
rect 511986 193058 512222 193294
rect 512306 193058 512542 193294
rect 511986 153378 512222 153614
rect 512306 153378 512542 153614
rect 511986 153058 512222 153294
rect 512306 153058 512542 153294
rect 511986 113378 512222 113614
rect 512306 113378 512542 113614
rect 511986 113058 512222 113294
rect 512306 113058 512542 113294
rect 511986 73378 512222 73614
rect 512306 73378 512542 73614
rect 511986 73058 512222 73294
rect 512306 73058 512542 73294
rect 511986 33378 512222 33614
rect 512306 33378 512542 33614
rect 511986 33058 512222 33294
rect 512306 33058 512542 33294
rect 491986 -6342 492222 -6106
rect 492306 -6342 492542 -6106
rect 491986 -6662 492222 -6426
rect 492306 -6662 492542 -6426
rect 520826 704602 521062 704838
rect 521146 704602 521382 704838
rect 520826 704282 521062 704518
rect 521146 704282 521382 704518
rect 520826 682218 521062 682454
rect 521146 682218 521382 682454
rect 520826 681898 521062 682134
rect 521146 681898 521382 682134
rect 520826 642218 521062 642454
rect 521146 642218 521382 642454
rect 520826 641898 521062 642134
rect 521146 641898 521382 642134
rect 520826 602218 521062 602454
rect 521146 602218 521382 602454
rect 520826 601898 521062 602134
rect 521146 601898 521382 602134
rect 520826 562218 521062 562454
rect 521146 562218 521382 562454
rect 520826 561898 521062 562134
rect 521146 561898 521382 562134
rect 520826 522218 521062 522454
rect 521146 522218 521382 522454
rect 520826 521898 521062 522134
rect 521146 521898 521382 522134
rect 520826 482218 521062 482454
rect 521146 482218 521382 482454
rect 520826 481898 521062 482134
rect 521146 481898 521382 482134
rect 520826 442218 521062 442454
rect 521146 442218 521382 442454
rect 520826 441898 521062 442134
rect 521146 441898 521382 442134
rect 520826 402218 521062 402454
rect 521146 402218 521382 402454
rect 520826 401898 521062 402134
rect 521146 401898 521382 402134
rect 520826 362218 521062 362454
rect 521146 362218 521382 362454
rect 520826 361898 521062 362134
rect 521146 361898 521382 362134
rect 520826 322218 521062 322454
rect 521146 322218 521382 322454
rect 520826 321898 521062 322134
rect 521146 321898 521382 322134
rect 520826 282218 521062 282454
rect 521146 282218 521382 282454
rect 520826 281898 521062 282134
rect 521146 281898 521382 282134
rect 520826 242218 521062 242454
rect 521146 242218 521382 242454
rect 520826 241898 521062 242134
rect 521146 241898 521382 242134
rect 520826 202218 521062 202454
rect 521146 202218 521382 202454
rect 520826 201898 521062 202134
rect 521146 201898 521382 202134
rect 520826 162218 521062 162454
rect 521146 162218 521382 162454
rect 520826 161898 521062 162134
rect 521146 161898 521382 162134
rect 520826 122218 521062 122454
rect 521146 122218 521382 122454
rect 520826 121898 521062 122134
rect 521146 121898 521382 122134
rect 520826 82218 521062 82454
rect 521146 82218 521382 82454
rect 520826 81898 521062 82134
rect 521146 81898 521382 82134
rect 520826 42218 521062 42454
rect 521146 42218 521382 42454
rect 520826 41898 521062 42134
rect 521146 41898 521382 42134
rect 520826 2218 521062 2454
rect 521146 2218 521382 2454
rect 520826 1898 521062 2134
rect 521146 1898 521382 2134
rect 520826 -582 521062 -346
rect 521146 -582 521382 -346
rect 520826 -902 521062 -666
rect 521146 -902 521382 -666
rect 524546 685938 524782 686174
rect 524866 685938 525102 686174
rect 524546 685618 524782 685854
rect 524866 685618 525102 685854
rect 524546 645938 524782 646174
rect 524866 645938 525102 646174
rect 524546 645618 524782 645854
rect 524866 645618 525102 645854
rect 524546 605938 524782 606174
rect 524866 605938 525102 606174
rect 524546 605618 524782 605854
rect 524866 605618 525102 605854
rect 524546 565938 524782 566174
rect 524866 565938 525102 566174
rect 524546 565618 524782 565854
rect 524866 565618 525102 565854
rect 524546 525938 524782 526174
rect 524866 525938 525102 526174
rect 524546 525618 524782 525854
rect 524866 525618 525102 525854
rect 524546 485938 524782 486174
rect 524866 485938 525102 486174
rect 524546 485618 524782 485854
rect 524866 485618 525102 485854
rect 524546 445938 524782 446174
rect 524866 445938 525102 446174
rect 524546 445618 524782 445854
rect 524866 445618 525102 445854
rect 524546 405938 524782 406174
rect 524866 405938 525102 406174
rect 524546 405618 524782 405854
rect 524866 405618 525102 405854
rect 524546 365938 524782 366174
rect 524866 365938 525102 366174
rect 524546 365618 524782 365854
rect 524866 365618 525102 365854
rect 524546 325938 524782 326174
rect 524866 325938 525102 326174
rect 524546 325618 524782 325854
rect 524866 325618 525102 325854
rect 524546 285938 524782 286174
rect 524866 285938 525102 286174
rect 524546 285618 524782 285854
rect 524866 285618 525102 285854
rect 524546 245938 524782 246174
rect 524866 245938 525102 246174
rect 524546 245618 524782 245854
rect 524866 245618 525102 245854
rect 524546 205938 524782 206174
rect 524866 205938 525102 206174
rect 524546 205618 524782 205854
rect 524866 205618 525102 205854
rect 524546 165938 524782 166174
rect 524866 165938 525102 166174
rect 524546 165618 524782 165854
rect 524866 165618 525102 165854
rect 524546 125938 524782 126174
rect 524866 125938 525102 126174
rect 524546 125618 524782 125854
rect 524866 125618 525102 125854
rect 524546 85938 524782 86174
rect 524866 85938 525102 86174
rect 524546 85618 524782 85854
rect 524866 85618 525102 85854
rect 524546 45938 524782 46174
rect 524866 45938 525102 46174
rect 524546 45618 524782 45854
rect 524866 45618 525102 45854
rect 524546 5938 524782 6174
rect 524866 5938 525102 6174
rect 524546 5618 524782 5854
rect 524866 5618 525102 5854
rect 524546 -2502 524782 -2266
rect 524866 -2502 525102 -2266
rect 524546 -2822 524782 -2586
rect 524866 -2822 525102 -2586
rect 528266 689658 528502 689894
rect 528586 689658 528822 689894
rect 528266 689338 528502 689574
rect 528586 689338 528822 689574
rect 528266 649658 528502 649894
rect 528586 649658 528822 649894
rect 528266 649338 528502 649574
rect 528586 649338 528822 649574
rect 528266 609658 528502 609894
rect 528586 609658 528822 609894
rect 528266 609338 528502 609574
rect 528586 609338 528822 609574
rect 528266 569658 528502 569894
rect 528586 569658 528822 569894
rect 528266 569338 528502 569574
rect 528586 569338 528822 569574
rect 528266 529658 528502 529894
rect 528586 529658 528822 529894
rect 528266 529338 528502 529574
rect 528586 529338 528822 529574
rect 528266 489658 528502 489894
rect 528586 489658 528822 489894
rect 528266 489338 528502 489574
rect 528586 489338 528822 489574
rect 528266 449658 528502 449894
rect 528586 449658 528822 449894
rect 528266 449338 528502 449574
rect 528586 449338 528822 449574
rect 528266 409658 528502 409894
rect 528586 409658 528822 409894
rect 528266 409338 528502 409574
rect 528586 409338 528822 409574
rect 528266 369658 528502 369894
rect 528586 369658 528822 369894
rect 528266 369338 528502 369574
rect 528586 369338 528822 369574
rect 528266 329658 528502 329894
rect 528586 329658 528822 329894
rect 528266 329338 528502 329574
rect 528586 329338 528822 329574
rect 528266 289658 528502 289894
rect 528586 289658 528822 289894
rect 528266 289338 528502 289574
rect 528586 289338 528822 289574
rect 528266 249658 528502 249894
rect 528586 249658 528822 249894
rect 528266 249338 528502 249574
rect 528586 249338 528822 249574
rect 528266 209658 528502 209894
rect 528586 209658 528822 209894
rect 528266 209338 528502 209574
rect 528586 209338 528822 209574
rect 528266 169658 528502 169894
rect 528586 169658 528822 169894
rect 528266 169338 528502 169574
rect 528586 169338 528822 169574
rect 528266 129658 528502 129894
rect 528586 129658 528822 129894
rect 528266 129338 528502 129574
rect 528586 129338 528822 129574
rect 528266 89658 528502 89894
rect 528586 89658 528822 89894
rect 528266 89338 528502 89574
rect 528586 89338 528822 89574
rect 528266 49658 528502 49894
rect 528586 49658 528822 49894
rect 528266 49338 528502 49574
rect 528586 49338 528822 49574
rect 528266 9658 528502 9894
rect 528586 9658 528822 9894
rect 528266 9338 528502 9574
rect 528586 9338 528822 9574
rect 528266 -4422 528502 -4186
rect 528586 -4422 528822 -4186
rect 528266 -4742 528502 -4506
rect 528586 -4742 528822 -4506
rect 551986 711322 552222 711558
rect 552306 711322 552542 711558
rect 551986 711002 552222 711238
rect 552306 711002 552542 711238
rect 548266 709402 548502 709638
rect 548586 709402 548822 709638
rect 548266 709082 548502 709318
rect 548586 709082 548822 709318
rect 544546 707482 544782 707718
rect 544866 707482 545102 707718
rect 544546 707162 544782 707398
rect 544866 707162 545102 707398
rect 531986 693378 532222 693614
rect 532306 693378 532542 693614
rect 531986 693058 532222 693294
rect 532306 693058 532542 693294
rect 531986 653378 532222 653614
rect 532306 653378 532542 653614
rect 531986 653058 532222 653294
rect 532306 653058 532542 653294
rect 531986 613378 532222 613614
rect 532306 613378 532542 613614
rect 531986 613058 532222 613294
rect 532306 613058 532542 613294
rect 531986 573378 532222 573614
rect 532306 573378 532542 573614
rect 531986 573058 532222 573294
rect 532306 573058 532542 573294
rect 531986 533378 532222 533614
rect 532306 533378 532542 533614
rect 531986 533058 532222 533294
rect 532306 533058 532542 533294
rect 531986 493378 532222 493614
rect 532306 493378 532542 493614
rect 531986 493058 532222 493294
rect 532306 493058 532542 493294
rect 531986 453378 532222 453614
rect 532306 453378 532542 453614
rect 531986 453058 532222 453294
rect 532306 453058 532542 453294
rect 531986 413378 532222 413614
rect 532306 413378 532542 413614
rect 531986 413058 532222 413294
rect 532306 413058 532542 413294
rect 531986 373378 532222 373614
rect 532306 373378 532542 373614
rect 531986 373058 532222 373294
rect 532306 373058 532542 373294
rect 531986 333378 532222 333614
rect 532306 333378 532542 333614
rect 531986 333058 532222 333294
rect 532306 333058 532542 333294
rect 531986 293378 532222 293614
rect 532306 293378 532542 293614
rect 531986 293058 532222 293294
rect 532306 293058 532542 293294
rect 531986 253378 532222 253614
rect 532306 253378 532542 253614
rect 531986 253058 532222 253294
rect 532306 253058 532542 253294
rect 531986 213378 532222 213614
rect 532306 213378 532542 213614
rect 531986 213058 532222 213294
rect 532306 213058 532542 213294
rect 531986 173378 532222 173614
rect 532306 173378 532542 173614
rect 531986 173058 532222 173294
rect 532306 173058 532542 173294
rect 531986 133378 532222 133614
rect 532306 133378 532542 133614
rect 531986 133058 532222 133294
rect 532306 133058 532542 133294
rect 531986 93378 532222 93614
rect 532306 93378 532542 93614
rect 531986 93058 532222 93294
rect 532306 93058 532542 93294
rect 531986 53378 532222 53614
rect 532306 53378 532542 53614
rect 531986 53058 532222 53294
rect 532306 53058 532542 53294
rect 531986 13378 532222 13614
rect 532306 13378 532542 13614
rect 531986 13058 532222 13294
rect 532306 13058 532542 13294
rect 511986 -7302 512222 -7066
rect 512306 -7302 512542 -7066
rect 511986 -7622 512222 -7386
rect 512306 -7622 512542 -7386
rect 540826 705562 541062 705798
rect 541146 705562 541382 705798
rect 540826 705242 541062 705478
rect 541146 705242 541382 705478
rect 540826 662218 541062 662454
rect 541146 662218 541382 662454
rect 540826 661898 541062 662134
rect 541146 661898 541382 662134
rect 540826 622218 541062 622454
rect 541146 622218 541382 622454
rect 540826 621898 541062 622134
rect 541146 621898 541382 622134
rect 540826 582218 541062 582454
rect 541146 582218 541382 582454
rect 540826 581898 541062 582134
rect 541146 581898 541382 582134
rect 540826 542218 541062 542454
rect 541146 542218 541382 542454
rect 540826 541898 541062 542134
rect 541146 541898 541382 542134
rect 540826 502218 541062 502454
rect 541146 502218 541382 502454
rect 540826 501898 541062 502134
rect 541146 501898 541382 502134
rect 540826 462218 541062 462454
rect 541146 462218 541382 462454
rect 540826 461898 541062 462134
rect 541146 461898 541382 462134
rect 540826 422218 541062 422454
rect 541146 422218 541382 422454
rect 540826 421898 541062 422134
rect 541146 421898 541382 422134
rect 540826 382218 541062 382454
rect 541146 382218 541382 382454
rect 540826 381898 541062 382134
rect 541146 381898 541382 382134
rect 540826 342218 541062 342454
rect 541146 342218 541382 342454
rect 540826 341898 541062 342134
rect 541146 341898 541382 342134
rect 540826 302218 541062 302454
rect 541146 302218 541382 302454
rect 540826 301898 541062 302134
rect 541146 301898 541382 302134
rect 540826 262218 541062 262454
rect 541146 262218 541382 262454
rect 540826 261898 541062 262134
rect 541146 261898 541382 262134
rect 540826 222218 541062 222454
rect 541146 222218 541382 222454
rect 540826 221898 541062 222134
rect 541146 221898 541382 222134
rect 540826 182218 541062 182454
rect 541146 182218 541382 182454
rect 540826 181898 541062 182134
rect 541146 181898 541382 182134
rect 540826 142218 541062 142454
rect 541146 142218 541382 142454
rect 540826 141898 541062 142134
rect 541146 141898 541382 142134
rect 540826 102218 541062 102454
rect 541146 102218 541382 102454
rect 540826 101898 541062 102134
rect 541146 101898 541382 102134
rect 540826 62218 541062 62454
rect 541146 62218 541382 62454
rect 540826 61898 541062 62134
rect 541146 61898 541382 62134
rect 540826 22218 541062 22454
rect 541146 22218 541382 22454
rect 540826 21898 541062 22134
rect 541146 21898 541382 22134
rect 540826 -1542 541062 -1306
rect 541146 -1542 541382 -1306
rect 540826 -1862 541062 -1626
rect 541146 -1862 541382 -1626
rect 544546 665938 544782 666174
rect 544866 665938 545102 666174
rect 544546 665618 544782 665854
rect 544866 665618 545102 665854
rect 544546 625938 544782 626174
rect 544866 625938 545102 626174
rect 544546 625618 544782 625854
rect 544866 625618 545102 625854
rect 544546 585938 544782 586174
rect 544866 585938 545102 586174
rect 544546 585618 544782 585854
rect 544866 585618 545102 585854
rect 544546 545938 544782 546174
rect 544866 545938 545102 546174
rect 544546 545618 544782 545854
rect 544866 545618 545102 545854
rect 544546 505938 544782 506174
rect 544866 505938 545102 506174
rect 544546 505618 544782 505854
rect 544866 505618 545102 505854
rect 544546 465938 544782 466174
rect 544866 465938 545102 466174
rect 544546 465618 544782 465854
rect 544866 465618 545102 465854
rect 544546 425938 544782 426174
rect 544866 425938 545102 426174
rect 544546 425618 544782 425854
rect 544866 425618 545102 425854
rect 544546 385938 544782 386174
rect 544866 385938 545102 386174
rect 544546 385618 544782 385854
rect 544866 385618 545102 385854
rect 544546 345938 544782 346174
rect 544866 345938 545102 346174
rect 544546 345618 544782 345854
rect 544866 345618 545102 345854
rect 544546 305938 544782 306174
rect 544866 305938 545102 306174
rect 544546 305618 544782 305854
rect 544866 305618 545102 305854
rect 544546 265938 544782 266174
rect 544866 265938 545102 266174
rect 544546 265618 544782 265854
rect 544866 265618 545102 265854
rect 544546 225938 544782 226174
rect 544866 225938 545102 226174
rect 544546 225618 544782 225854
rect 544866 225618 545102 225854
rect 544546 185938 544782 186174
rect 544866 185938 545102 186174
rect 544546 185618 544782 185854
rect 544866 185618 545102 185854
rect 544546 145938 544782 146174
rect 544866 145938 545102 146174
rect 544546 145618 544782 145854
rect 544866 145618 545102 145854
rect 544546 105938 544782 106174
rect 544866 105938 545102 106174
rect 544546 105618 544782 105854
rect 544866 105618 545102 105854
rect 544546 65938 544782 66174
rect 544866 65938 545102 66174
rect 544546 65618 544782 65854
rect 544866 65618 545102 65854
rect 544546 25938 544782 26174
rect 544866 25938 545102 26174
rect 544546 25618 544782 25854
rect 544866 25618 545102 25854
rect 544546 -3462 544782 -3226
rect 544866 -3462 545102 -3226
rect 544546 -3782 544782 -3546
rect 544866 -3782 545102 -3546
rect 548266 669658 548502 669894
rect 548586 669658 548822 669894
rect 548266 669338 548502 669574
rect 548586 669338 548822 669574
rect 548266 629658 548502 629894
rect 548586 629658 548822 629894
rect 548266 629338 548502 629574
rect 548586 629338 548822 629574
rect 548266 589658 548502 589894
rect 548586 589658 548822 589894
rect 548266 589338 548502 589574
rect 548586 589338 548822 589574
rect 548266 549658 548502 549894
rect 548586 549658 548822 549894
rect 548266 549338 548502 549574
rect 548586 549338 548822 549574
rect 548266 509658 548502 509894
rect 548586 509658 548822 509894
rect 548266 509338 548502 509574
rect 548586 509338 548822 509574
rect 548266 469658 548502 469894
rect 548586 469658 548822 469894
rect 548266 469338 548502 469574
rect 548586 469338 548822 469574
rect 548266 429658 548502 429894
rect 548586 429658 548822 429894
rect 548266 429338 548502 429574
rect 548586 429338 548822 429574
rect 548266 389658 548502 389894
rect 548586 389658 548822 389894
rect 548266 389338 548502 389574
rect 548586 389338 548822 389574
rect 548266 349658 548502 349894
rect 548586 349658 548822 349894
rect 548266 349338 548502 349574
rect 548586 349338 548822 349574
rect 548266 309658 548502 309894
rect 548586 309658 548822 309894
rect 548266 309338 548502 309574
rect 548586 309338 548822 309574
rect 548266 269658 548502 269894
rect 548586 269658 548822 269894
rect 548266 269338 548502 269574
rect 548586 269338 548822 269574
rect 548266 229658 548502 229894
rect 548586 229658 548822 229894
rect 548266 229338 548502 229574
rect 548586 229338 548822 229574
rect 548266 189658 548502 189894
rect 548586 189658 548822 189894
rect 548266 189338 548502 189574
rect 548586 189338 548822 189574
rect 548266 149658 548502 149894
rect 548586 149658 548822 149894
rect 548266 149338 548502 149574
rect 548586 149338 548822 149574
rect 548266 109658 548502 109894
rect 548586 109658 548822 109894
rect 548266 109338 548502 109574
rect 548586 109338 548822 109574
rect 548266 69658 548502 69894
rect 548586 69658 548822 69894
rect 548266 69338 548502 69574
rect 548586 69338 548822 69574
rect 548266 29658 548502 29894
rect 548586 29658 548822 29894
rect 548266 29338 548502 29574
rect 548586 29338 548822 29574
rect 548266 -5382 548502 -5146
rect 548586 -5382 548822 -5146
rect 548266 -5702 548502 -5466
rect 548586 -5702 548822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 571986 710362 572222 710598
rect 572306 710362 572542 710598
rect 571986 710042 572222 710278
rect 572306 710042 572542 710278
rect 568266 708442 568502 708678
rect 568586 708442 568822 708678
rect 568266 708122 568502 708358
rect 568586 708122 568822 708358
rect 564546 706522 564782 706758
rect 564866 706522 565102 706758
rect 564546 706202 564782 706438
rect 564866 706202 565102 706438
rect 551986 673378 552222 673614
rect 552306 673378 552542 673614
rect 551986 673058 552222 673294
rect 552306 673058 552542 673294
rect 551986 633378 552222 633614
rect 552306 633378 552542 633614
rect 551986 633058 552222 633294
rect 552306 633058 552542 633294
rect 551986 593378 552222 593614
rect 552306 593378 552542 593614
rect 551986 593058 552222 593294
rect 552306 593058 552542 593294
rect 551986 553378 552222 553614
rect 552306 553378 552542 553614
rect 551986 553058 552222 553294
rect 552306 553058 552542 553294
rect 551986 513378 552222 513614
rect 552306 513378 552542 513614
rect 551986 513058 552222 513294
rect 552306 513058 552542 513294
rect 551986 473378 552222 473614
rect 552306 473378 552542 473614
rect 551986 473058 552222 473294
rect 552306 473058 552542 473294
rect 551986 433378 552222 433614
rect 552306 433378 552542 433614
rect 551986 433058 552222 433294
rect 552306 433058 552542 433294
rect 551986 393378 552222 393614
rect 552306 393378 552542 393614
rect 551986 393058 552222 393294
rect 552306 393058 552542 393294
rect 551986 353378 552222 353614
rect 552306 353378 552542 353614
rect 551986 353058 552222 353294
rect 552306 353058 552542 353294
rect 551986 313378 552222 313614
rect 552306 313378 552542 313614
rect 551986 313058 552222 313294
rect 552306 313058 552542 313294
rect 551986 273378 552222 273614
rect 552306 273378 552542 273614
rect 551986 273058 552222 273294
rect 552306 273058 552542 273294
rect 551986 233378 552222 233614
rect 552306 233378 552542 233614
rect 551986 233058 552222 233294
rect 552306 233058 552542 233294
rect 551986 193378 552222 193614
rect 552306 193378 552542 193614
rect 551986 193058 552222 193294
rect 552306 193058 552542 193294
rect 551986 153378 552222 153614
rect 552306 153378 552542 153614
rect 551986 153058 552222 153294
rect 552306 153058 552542 153294
rect 551986 113378 552222 113614
rect 552306 113378 552542 113614
rect 551986 113058 552222 113294
rect 552306 113058 552542 113294
rect 551986 73378 552222 73614
rect 552306 73378 552542 73614
rect 551986 73058 552222 73294
rect 552306 73058 552542 73294
rect 551986 33378 552222 33614
rect 552306 33378 552542 33614
rect 551986 33058 552222 33294
rect 552306 33058 552542 33294
rect 531986 -6342 532222 -6106
rect 532306 -6342 532542 -6106
rect 531986 -6662 532222 -6426
rect 532306 -6662 532542 -6426
rect 560826 704602 561062 704838
rect 561146 704602 561382 704838
rect 560826 704282 561062 704518
rect 561146 704282 561382 704518
rect 560826 682218 561062 682454
rect 561146 682218 561382 682454
rect 560826 681898 561062 682134
rect 561146 681898 561382 682134
rect 560826 642218 561062 642454
rect 561146 642218 561382 642454
rect 560826 641898 561062 642134
rect 561146 641898 561382 642134
rect 560826 602218 561062 602454
rect 561146 602218 561382 602454
rect 560826 601898 561062 602134
rect 561146 601898 561382 602134
rect 560826 562218 561062 562454
rect 561146 562218 561382 562454
rect 560826 561898 561062 562134
rect 561146 561898 561382 562134
rect 560826 522218 561062 522454
rect 561146 522218 561382 522454
rect 560826 521898 561062 522134
rect 561146 521898 561382 522134
rect 560826 482218 561062 482454
rect 561146 482218 561382 482454
rect 560826 481898 561062 482134
rect 561146 481898 561382 482134
rect 560826 442218 561062 442454
rect 561146 442218 561382 442454
rect 560826 441898 561062 442134
rect 561146 441898 561382 442134
rect 560826 402218 561062 402454
rect 561146 402218 561382 402454
rect 560826 401898 561062 402134
rect 561146 401898 561382 402134
rect 560826 362218 561062 362454
rect 561146 362218 561382 362454
rect 560826 361898 561062 362134
rect 561146 361898 561382 362134
rect 560826 322218 561062 322454
rect 561146 322218 561382 322454
rect 560826 321898 561062 322134
rect 561146 321898 561382 322134
rect 560826 282218 561062 282454
rect 561146 282218 561382 282454
rect 560826 281898 561062 282134
rect 561146 281898 561382 282134
rect 560826 242218 561062 242454
rect 561146 242218 561382 242454
rect 560826 241898 561062 242134
rect 561146 241898 561382 242134
rect 560826 202218 561062 202454
rect 561146 202218 561382 202454
rect 560826 201898 561062 202134
rect 561146 201898 561382 202134
rect 560826 162218 561062 162454
rect 561146 162218 561382 162454
rect 560826 161898 561062 162134
rect 561146 161898 561382 162134
rect 560826 122218 561062 122454
rect 561146 122218 561382 122454
rect 560826 121898 561062 122134
rect 561146 121898 561382 122134
rect 560826 82218 561062 82454
rect 561146 82218 561382 82454
rect 560826 81898 561062 82134
rect 561146 81898 561382 82134
rect 560826 42218 561062 42454
rect 561146 42218 561382 42454
rect 560826 41898 561062 42134
rect 561146 41898 561382 42134
rect 560826 2218 561062 2454
rect 561146 2218 561382 2454
rect 560826 1898 561062 2134
rect 561146 1898 561382 2134
rect 560826 -582 561062 -346
rect 561146 -582 561382 -346
rect 560826 -902 561062 -666
rect 561146 -902 561382 -666
rect 564546 685938 564782 686174
rect 564866 685938 565102 686174
rect 564546 685618 564782 685854
rect 564866 685618 565102 685854
rect 564546 645938 564782 646174
rect 564866 645938 565102 646174
rect 564546 645618 564782 645854
rect 564866 645618 565102 645854
rect 564546 605938 564782 606174
rect 564866 605938 565102 606174
rect 564546 605618 564782 605854
rect 564866 605618 565102 605854
rect 564546 565938 564782 566174
rect 564866 565938 565102 566174
rect 564546 565618 564782 565854
rect 564866 565618 565102 565854
rect 564546 525938 564782 526174
rect 564866 525938 565102 526174
rect 564546 525618 564782 525854
rect 564866 525618 565102 525854
rect 564546 485938 564782 486174
rect 564866 485938 565102 486174
rect 564546 485618 564782 485854
rect 564866 485618 565102 485854
rect 564546 445938 564782 446174
rect 564866 445938 565102 446174
rect 564546 445618 564782 445854
rect 564866 445618 565102 445854
rect 564546 405938 564782 406174
rect 564866 405938 565102 406174
rect 564546 405618 564782 405854
rect 564866 405618 565102 405854
rect 564546 365938 564782 366174
rect 564866 365938 565102 366174
rect 564546 365618 564782 365854
rect 564866 365618 565102 365854
rect 564546 325938 564782 326174
rect 564866 325938 565102 326174
rect 564546 325618 564782 325854
rect 564866 325618 565102 325854
rect 564546 285938 564782 286174
rect 564866 285938 565102 286174
rect 564546 285618 564782 285854
rect 564866 285618 565102 285854
rect 564546 245938 564782 246174
rect 564866 245938 565102 246174
rect 564546 245618 564782 245854
rect 564866 245618 565102 245854
rect 564546 205938 564782 206174
rect 564866 205938 565102 206174
rect 564546 205618 564782 205854
rect 564866 205618 565102 205854
rect 564546 165938 564782 166174
rect 564866 165938 565102 166174
rect 564546 165618 564782 165854
rect 564866 165618 565102 165854
rect 564546 125938 564782 126174
rect 564866 125938 565102 126174
rect 564546 125618 564782 125854
rect 564866 125618 565102 125854
rect 564546 85938 564782 86174
rect 564866 85938 565102 86174
rect 564546 85618 564782 85854
rect 564866 85618 565102 85854
rect 564546 45938 564782 46174
rect 564866 45938 565102 46174
rect 564546 45618 564782 45854
rect 564866 45618 565102 45854
rect 564546 5938 564782 6174
rect 564866 5938 565102 6174
rect 564546 5618 564782 5854
rect 564866 5618 565102 5854
rect 564546 -2502 564782 -2266
rect 564866 -2502 565102 -2266
rect 564546 -2822 564782 -2586
rect 564866 -2822 565102 -2586
rect 568266 689658 568502 689894
rect 568586 689658 568822 689894
rect 568266 689338 568502 689574
rect 568586 689338 568822 689574
rect 568266 649658 568502 649894
rect 568586 649658 568822 649894
rect 568266 649338 568502 649574
rect 568586 649338 568822 649574
rect 568266 609658 568502 609894
rect 568586 609658 568822 609894
rect 568266 609338 568502 609574
rect 568586 609338 568822 609574
rect 568266 569658 568502 569894
rect 568586 569658 568822 569894
rect 568266 569338 568502 569574
rect 568586 569338 568822 569574
rect 568266 529658 568502 529894
rect 568586 529658 568822 529894
rect 568266 529338 568502 529574
rect 568586 529338 568822 529574
rect 568266 489658 568502 489894
rect 568586 489658 568822 489894
rect 568266 489338 568502 489574
rect 568586 489338 568822 489574
rect 568266 449658 568502 449894
rect 568586 449658 568822 449894
rect 568266 449338 568502 449574
rect 568586 449338 568822 449574
rect 568266 409658 568502 409894
rect 568586 409658 568822 409894
rect 568266 409338 568502 409574
rect 568586 409338 568822 409574
rect 568266 369658 568502 369894
rect 568586 369658 568822 369894
rect 568266 369338 568502 369574
rect 568586 369338 568822 369574
rect 568266 329658 568502 329894
rect 568586 329658 568822 329894
rect 568266 329338 568502 329574
rect 568586 329338 568822 329574
rect 568266 289658 568502 289894
rect 568586 289658 568822 289894
rect 568266 289338 568502 289574
rect 568586 289338 568822 289574
rect 568266 249658 568502 249894
rect 568586 249658 568822 249894
rect 568266 249338 568502 249574
rect 568586 249338 568822 249574
rect 568266 209658 568502 209894
rect 568586 209658 568822 209894
rect 568266 209338 568502 209574
rect 568586 209338 568822 209574
rect 568266 169658 568502 169894
rect 568586 169658 568822 169894
rect 568266 169338 568502 169574
rect 568586 169338 568822 169574
rect 568266 129658 568502 129894
rect 568586 129658 568822 129894
rect 568266 129338 568502 129574
rect 568586 129338 568822 129574
rect 568266 89658 568502 89894
rect 568586 89658 568822 89894
rect 568266 89338 568502 89574
rect 568586 89338 568822 89574
rect 568266 49658 568502 49894
rect 568586 49658 568822 49894
rect 568266 49338 568502 49574
rect 568586 49338 568822 49574
rect 568266 9658 568502 9894
rect 568586 9658 568822 9894
rect 568266 9338 568502 9574
rect 568586 9338 568822 9574
rect 568266 -4422 568502 -4186
rect 568586 -4422 568822 -4186
rect 568266 -4742 568502 -4506
rect 568586 -4742 568822 -4506
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 571986 693378 572222 693614
rect 572306 693378 572542 693614
rect 571986 693058 572222 693294
rect 572306 693058 572542 693294
rect 571986 653378 572222 653614
rect 572306 653378 572542 653614
rect 571986 653058 572222 653294
rect 572306 653058 572542 653294
rect 571986 613378 572222 613614
rect 572306 613378 572542 613614
rect 571986 613058 572222 613294
rect 572306 613058 572542 613294
rect 571986 573378 572222 573614
rect 572306 573378 572542 573614
rect 571986 573058 572222 573294
rect 572306 573058 572542 573294
rect 571986 533378 572222 533614
rect 572306 533378 572542 533614
rect 571986 533058 572222 533294
rect 572306 533058 572542 533294
rect 571986 493378 572222 493614
rect 572306 493378 572542 493614
rect 571986 493058 572222 493294
rect 572306 493058 572542 493294
rect 571986 453378 572222 453614
rect 572306 453378 572542 453614
rect 571986 453058 572222 453294
rect 572306 453058 572542 453294
rect 571986 413378 572222 413614
rect 572306 413378 572542 413614
rect 571986 413058 572222 413294
rect 572306 413058 572542 413294
rect 571986 373378 572222 373614
rect 572306 373378 572542 373614
rect 571986 373058 572222 373294
rect 572306 373058 572542 373294
rect 571986 333378 572222 333614
rect 572306 333378 572542 333614
rect 571986 333058 572222 333294
rect 572306 333058 572542 333294
rect 571986 293378 572222 293614
rect 572306 293378 572542 293614
rect 571986 293058 572222 293294
rect 572306 293058 572542 293294
rect 571986 253378 572222 253614
rect 572306 253378 572542 253614
rect 571986 253058 572222 253294
rect 572306 253058 572542 253294
rect 571986 213378 572222 213614
rect 572306 213378 572542 213614
rect 571986 213058 572222 213294
rect 572306 213058 572542 213294
rect 571986 173378 572222 173614
rect 572306 173378 572542 173614
rect 571986 173058 572222 173294
rect 572306 173058 572542 173294
rect 571986 133378 572222 133614
rect 572306 133378 572542 133614
rect 571986 133058 572222 133294
rect 572306 133058 572542 133294
rect 571986 93378 572222 93614
rect 572306 93378 572542 93614
rect 571986 93058 572222 93294
rect 572306 93058 572542 93294
rect 571986 53378 572222 53614
rect 572306 53378 572542 53614
rect 571986 53058 572222 53294
rect 572306 53058 572542 53294
rect 571986 13378 572222 13614
rect 572306 13378 572542 13614
rect 571986 13058 572222 13294
rect 572306 13058 572542 13294
rect 551986 -7302 552222 -7066
rect 552306 -7302 552542 -7066
rect 551986 -7622 552222 -7386
rect 552306 -7622 552542 -7386
rect 580826 705562 581062 705798
rect 581146 705562 581382 705798
rect 580826 705242 581062 705478
rect 581146 705242 581382 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 580826 662218 581062 662454
rect 581146 662218 581382 662454
rect 580826 661898 581062 662134
rect 581146 661898 581382 662134
rect 580826 622218 581062 622454
rect 581146 622218 581382 622454
rect 580826 621898 581062 622134
rect 581146 621898 581382 622134
rect 580826 582218 581062 582454
rect 581146 582218 581382 582454
rect 580826 581898 581062 582134
rect 581146 581898 581382 582134
rect 580826 542218 581062 542454
rect 581146 542218 581382 542454
rect 580826 541898 581062 542134
rect 581146 541898 581382 542134
rect 580826 502218 581062 502454
rect 581146 502218 581382 502454
rect 580826 501898 581062 502134
rect 581146 501898 581382 502134
rect 580826 462218 581062 462454
rect 581146 462218 581382 462454
rect 580826 461898 581062 462134
rect 581146 461898 581382 462134
rect 580826 422218 581062 422454
rect 581146 422218 581382 422454
rect 580826 421898 581062 422134
rect 581146 421898 581382 422134
rect 580826 382218 581062 382454
rect 581146 382218 581382 382454
rect 580826 381898 581062 382134
rect 581146 381898 581382 382134
rect 580826 342218 581062 342454
rect 581146 342218 581382 342454
rect 580826 341898 581062 342134
rect 581146 341898 581382 342134
rect 580826 302218 581062 302454
rect 581146 302218 581382 302454
rect 580826 301898 581062 302134
rect 581146 301898 581382 302134
rect 580826 262218 581062 262454
rect 581146 262218 581382 262454
rect 580826 261898 581062 262134
rect 581146 261898 581382 262134
rect 580826 222218 581062 222454
rect 581146 222218 581382 222454
rect 580826 221898 581062 222134
rect 581146 221898 581382 222134
rect 580826 182218 581062 182454
rect 581146 182218 581382 182454
rect 580826 181898 581062 182134
rect 581146 181898 581382 182134
rect 580826 142218 581062 142454
rect 581146 142218 581382 142454
rect 580826 141898 581062 142134
rect 581146 141898 581382 142134
rect 580826 102218 581062 102454
rect 581146 102218 581382 102454
rect 580826 101898 581062 102134
rect 581146 101898 581382 102134
rect 580826 62218 581062 62454
rect 581146 62218 581382 62454
rect 580826 61898 581062 62134
rect 581146 61898 581382 62134
rect 580826 22218 581062 22454
rect 581146 22218 581382 22454
rect 580826 21898 581062 22134
rect 581146 21898 581382 22134
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 682218 585578 682454
rect 585662 682218 585898 682454
rect 585342 681898 585578 682134
rect 585662 681898 585898 682134
rect 585342 642218 585578 642454
rect 585662 642218 585898 642454
rect 585342 641898 585578 642134
rect 585662 641898 585898 642134
rect 585342 602218 585578 602454
rect 585662 602218 585898 602454
rect 585342 601898 585578 602134
rect 585662 601898 585898 602134
rect 585342 562218 585578 562454
rect 585662 562218 585898 562454
rect 585342 561898 585578 562134
rect 585662 561898 585898 562134
rect 585342 522218 585578 522454
rect 585662 522218 585898 522454
rect 585342 521898 585578 522134
rect 585662 521898 585898 522134
rect 585342 482218 585578 482454
rect 585662 482218 585898 482454
rect 585342 481898 585578 482134
rect 585662 481898 585898 482134
rect 585342 442218 585578 442454
rect 585662 442218 585898 442454
rect 585342 441898 585578 442134
rect 585662 441898 585898 442134
rect 585342 402218 585578 402454
rect 585662 402218 585898 402454
rect 585342 401898 585578 402134
rect 585662 401898 585898 402134
rect 585342 362218 585578 362454
rect 585662 362218 585898 362454
rect 585342 361898 585578 362134
rect 585662 361898 585898 362134
rect 585342 322218 585578 322454
rect 585662 322218 585898 322454
rect 585342 321898 585578 322134
rect 585662 321898 585898 322134
rect 585342 282218 585578 282454
rect 585662 282218 585898 282454
rect 585342 281898 585578 282134
rect 585662 281898 585898 282134
rect 585342 242218 585578 242454
rect 585662 242218 585898 242454
rect 585342 241898 585578 242134
rect 585662 241898 585898 242134
rect 585342 202218 585578 202454
rect 585662 202218 585898 202454
rect 585342 201898 585578 202134
rect 585662 201898 585898 202134
rect 585342 162218 585578 162454
rect 585662 162218 585898 162454
rect 585342 161898 585578 162134
rect 585662 161898 585898 162134
rect 585342 122218 585578 122454
rect 585662 122218 585898 122454
rect 585342 121898 585578 122134
rect 585662 121898 585898 122134
rect 585342 82218 585578 82454
rect 585662 82218 585898 82454
rect 585342 81898 585578 82134
rect 585662 81898 585898 82134
rect 585342 42218 585578 42454
rect 585662 42218 585898 42454
rect 585342 41898 585578 42134
rect 585662 41898 585898 42134
rect 585342 2218 585578 2454
rect 585662 2218 585898 2454
rect 585342 1898 585578 2134
rect 585662 1898 585898 2134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 662218 586538 662454
rect 586622 662218 586858 662454
rect 586302 661898 586538 662134
rect 586622 661898 586858 662134
rect 586302 622218 586538 622454
rect 586622 622218 586858 622454
rect 586302 621898 586538 622134
rect 586622 621898 586858 622134
rect 586302 582218 586538 582454
rect 586622 582218 586858 582454
rect 586302 581898 586538 582134
rect 586622 581898 586858 582134
rect 586302 542218 586538 542454
rect 586622 542218 586858 542454
rect 586302 541898 586538 542134
rect 586622 541898 586858 542134
rect 586302 502218 586538 502454
rect 586622 502218 586858 502454
rect 586302 501898 586538 502134
rect 586622 501898 586858 502134
rect 586302 462218 586538 462454
rect 586622 462218 586858 462454
rect 586302 461898 586538 462134
rect 586622 461898 586858 462134
rect 586302 422218 586538 422454
rect 586622 422218 586858 422454
rect 586302 421898 586538 422134
rect 586622 421898 586858 422134
rect 586302 382218 586538 382454
rect 586622 382218 586858 382454
rect 586302 381898 586538 382134
rect 586622 381898 586858 382134
rect 586302 342218 586538 342454
rect 586622 342218 586858 342454
rect 586302 341898 586538 342134
rect 586622 341898 586858 342134
rect 586302 302218 586538 302454
rect 586622 302218 586858 302454
rect 586302 301898 586538 302134
rect 586622 301898 586858 302134
rect 586302 262218 586538 262454
rect 586622 262218 586858 262454
rect 586302 261898 586538 262134
rect 586622 261898 586858 262134
rect 586302 222218 586538 222454
rect 586622 222218 586858 222454
rect 586302 221898 586538 222134
rect 586622 221898 586858 222134
rect 586302 182218 586538 182454
rect 586622 182218 586858 182454
rect 586302 181898 586538 182134
rect 586622 181898 586858 182134
rect 586302 142218 586538 142454
rect 586622 142218 586858 142454
rect 586302 141898 586538 142134
rect 586622 141898 586858 142134
rect 586302 102218 586538 102454
rect 586622 102218 586858 102454
rect 586302 101898 586538 102134
rect 586622 101898 586858 102134
rect 586302 62218 586538 62454
rect 586622 62218 586858 62454
rect 586302 61898 586538 62134
rect 586622 61898 586858 62134
rect 586302 22218 586538 22454
rect 586622 22218 586858 22454
rect 586302 21898 586538 22134
rect 586622 21898 586858 22134
rect 580826 -1542 581062 -1306
rect 581146 -1542 581382 -1306
rect 580826 -1862 581062 -1626
rect 581146 -1862 581382 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 685938 587498 686174
rect 587582 685938 587818 686174
rect 587262 685618 587498 685854
rect 587582 685618 587818 685854
rect 587262 645938 587498 646174
rect 587582 645938 587818 646174
rect 587262 645618 587498 645854
rect 587582 645618 587818 645854
rect 587262 605938 587498 606174
rect 587582 605938 587818 606174
rect 587262 605618 587498 605854
rect 587582 605618 587818 605854
rect 587262 565938 587498 566174
rect 587582 565938 587818 566174
rect 587262 565618 587498 565854
rect 587582 565618 587818 565854
rect 587262 525938 587498 526174
rect 587582 525938 587818 526174
rect 587262 525618 587498 525854
rect 587582 525618 587818 525854
rect 587262 485938 587498 486174
rect 587582 485938 587818 486174
rect 587262 485618 587498 485854
rect 587582 485618 587818 485854
rect 587262 445938 587498 446174
rect 587582 445938 587818 446174
rect 587262 445618 587498 445854
rect 587582 445618 587818 445854
rect 587262 405938 587498 406174
rect 587582 405938 587818 406174
rect 587262 405618 587498 405854
rect 587582 405618 587818 405854
rect 587262 365938 587498 366174
rect 587582 365938 587818 366174
rect 587262 365618 587498 365854
rect 587582 365618 587818 365854
rect 587262 325938 587498 326174
rect 587582 325938 587818 326174
rect 587262 325618 587498 325854
rect 587582 325618 587818 325854
rect 587262 285938 587498 286174
rect 587582 285938 587818 286174
rect 587262 285618 587498 285854
rect 587582 285618 587818 285854
rect 587262 245938 587498 246174
rect 587582 245938 587818 246174
rect 587262 245618 587498 245854
rect 587582 245618 587818 245854
rect 587262 205938 587498 206174
rect 587582 205938 587818 206174
rect 587262 205618 587498 205854
rect 587582 205618 587818 205854
rect 587262 165938 587498 166174
rect 587582 165938 587818 166174
rect 587262 165618 587498 165854
rect 587582 165618 587818 165854
rect 587262 125938 587498 126174
rect 587582 125938 587818 126174
rect 587262 125618 587498 125854
rect 587582 125618 587818 125854
rect 587262 85938 587498 86174
rect 587582 85938 587818 86174
rect 587262 85618 587498 85854
rect 587582 85618 587818 85854
rect 587262 45938 587498 46174
rect 587582 45938 587818 46174
rect 587262 45618 587498 45854
rect 587582 45618 587818 45854
rect 587262 5938 587498 6174
rect 587582 5938 587818 6174
rect 587262 5618 587498 5854
rect 587582 5618 587818 5854
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 665938 588458 666174
rect 588542 665938 588778 666174
rect 588222 665618 588458 665854
rect 588542 665618 588778 665854
rect 588222 625938 588458 626174
rect 588542 625938 588778 626174
rect 588222 625618 588458 625854
rect 588542 625618 588778 625854
rect 588222 585938 588458 586174
rect 588542 585938 588778 586174
rect 588222 585618 588458 585854
rect 588542 585618 588778 585854
rect 588222 545938 588458 546174
rect 588542 545938 588778 546174
rect 588222 545618 588458 545854
rect 588542 545618 588778 545854
rect 588222 505938 588458 506174
rect 588542 505938 588778 506174
rect 588222 505618 588458 505854
rect 588542 505618 588778 505854
rect 588222 465938 588458 466174
rect 588542 465938 588778 466174
rect 588222 465618 588458 465854
rect 588542 465618 588778 465854
rect 588222 425938 588458 426174
rect 588542 425938 588778 426174
rect 588222 425618 588458 425854
rect 588542 425618 588778 425854
rect 588222 385938 588458 386174
rect 588542 385938 588778 386174
rect 588222 385618 588458 385854
rect 588542 385618 588778 385854
rect 588222 345938 588458 346174
rect 588542 345938 588778 346174
rect 588222 345618 588458 345854
rect 588542 345618 588778 345854
rect 588222 305938 588458 306174
rect 588542 305938 588778 306174
rect 588222 305618 588458 305854
rect 588542 305618 588778 305854
rect 588222 265938 588458 266174
rect 588542 265938 588778 266174
rect 588222 265618 588458 265854
rect 588542 265618 588778 265854
rect 588222 225938 588458 226174
rect 588542 225938 588778 226174
rect 588222 225618 588458 225854
rect 588542 225618 588778 225854
rect 588222 185938 588458 186174
rect 588542 185938 588778 186174
rect 588222 185618 588458 185854
rect 588542 185618 588778 185854
rect 588222 145938 588458 146174
rect 588542 145938 588778 146174
rect 588222 145618 588458 145854
rect 588542 145618 588778 145854
rect 588222 105938 588458 106174
rect 588542 105938 588778 106174
rect 588222 105618 588458 105854
rect 588542 105618 588778 105854
rect 588222 65938 588458 66174
rect 588542 65938 588778 66174
rect 588222 65618 588458 65854
rect 588542 65618 588778 65854
rect 588222 25938 588458 26174
rect 588542 25938 588778 26174
rect 588222 25618 588458 25854
rect 588542 25618 588778 25854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 689658 589418 689894
rect 589502 689658 589738 689894
rect 589182 689338 589418 689574
rect 589502 689338 589738 689574
rect 589182 649658 589418 649894
rect 589502 649658 589738 649894
rect 589182 649338 589418 649574
rect 589502 649338 589738 649574
rect 589182 609658 589418 609894
rect 589502 609658 589738 609894
rect 589182 609338 589418 609574
rect 589502 609338 589738 609574
rect 589182 569658 589418 569894
rect 589502 569658 589738 569894
rect 589182 569338 589418 569574
rect 589502 569338 589738 569574
rect 589182 529658 589418 529894
rect 589502 529658 589738 529894
rect 589182 529338 589418 529574
rect 589502 529338 589738 529574
rect 589182 489658 589418 489894
rect 589502 489658 589738 489894
rect 589182 489338 589418 489574
rect 589502 489338 589738 489574
rect 589182 449658 589418 449894
rect 589502 449658 589738 449894
rect 589182 449338 589418 449574
rect 589502 449338 589738 449574
rect 589182 409658 589418 409894
rect 589502 409658 589738 409894
rect 589182 409338 589418 409574
rect 589502 409338 589738 409574
rect 589182 369658 589418 369894
rect 589502 369658 589738 369894
rect 589182 369338 589418 369574
rect 589502 369338 589738 369574
rect 589182 329658 589418 329894
rect 589502 329658 589738 329894
rect 589182 329338 589418 329574
rect 589502 329338 589738 329574
rect 589182 289658 589418 289894
rect 589502 289658 589738 289894
rect 589182 289338 589418 289574
rect 589502 289338 589738 289574
rect 589182 249658 589418 249894
rect 589502 249658 589738 249894
rect 589182 249338 589418 249574
rect 589502 249338 589738 249574
rect 589182 209658 589418 209894
rect 589502 209658 589738 209894
rect 589182 209338 589418 209574
rect 589502 209338 589738 209574
rect 589182 169658 589418 169894
rect 589502 169658 589738 169894
rect 589182 169338 589418 169574
rect 589502 169338 589738 169574
rect 589182 129658 589418 129894
rect 589502 129658 589738 129894
rect 589182 129338 589418 129574
rect 589502 129338 589738 129574
rect 589182 89658 589418 89894
rect 589502 89658 589738 89894
rect 589182 89338 589418 89574
rect 589502 89338 589738 89574
rect 589182 49658 589418 49894
rect 589502 49658 589738 49894
rect 589182 49338 589418 49574
rect 589502 49338 589738 49574
rect 589182 9658 589418 9894
rect 589502 9658 589738 9894
rect 589182 9338 589418 9574
rect 589502 9338 589738 9574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669658 590378 669894
rect 590462 669658 590698 669894
rect 590142 669338 590378 669574
rect 590462 669338 590698 669574
rect 590142 629658 590378 629894
rect 590462 629658 590698 629894
rect 590142 629338 590378 629574
rect 590462 629338 590698 629574
rect 590142 589658 590378 589894
rect 590462 589658 590698 589894
rect 590142 589338 590378 589574
rect 590462 589338 590698 589574
rect 590142 549658 590378 549894
rect 590462 549658 590698 549894
rect 590142 549338 590378 549574
rect 590462 549338 590698 549574
rect 590142 509658 590378 509894
rect 590462 509658 590698 509894
rect 590142 509338 590378 509574
rect 590462 509338 590698 509574
rect 590142 469658 590378 469894
rect 590462 469658 590698 469894
rect 590142 469338 590378 469574
rect 590462 469338 590698 469574
rect 590142 429658 590378 429894
rect 590462 429658 590698 429894
rect 590142 429338 590378 429574
rect 590462 429338 590698 429574
rect 590142 389658 590378 389894
rect 590462 389658 590698 389894
rect 590142 389338 590378 389574
rect 590462 389338 590698 389574
rect 590142 349658 590378 349894
rect 590462 349658 590698 349894
rect 590142 349338 590378 349574
rect 590462 349338 590698 349574
rect 590142 309658 590378 309894
rect 590462 309658 590698 309894
rect 590142 309338 590378 309574
rect 590462 309338 590698 309574
rect 590142 269658 590378 269894
rect 590462 269658 590698 269894
rect 590142 269338 590378 269574
rect 590462 269338 590698 269574
rect 590142 229658 590378 229894
rect 590462 229658 590698 229894
rect 590142 229338 590378 229574
rect 590462 229338 590698 229574
rect 590142 189658 590378 189894
rect 590462 189658 590698 189894
rect 590142 189338 590378 189574
rect 590462 189338 590698 189574
rect 590142 149658 590378 149894
rect 590462 149658 590698 149894
rect 590142 149338 590378 149574
rect 590462 149338 590698 149574
rect 590142 109658 590378 109894
rect 590462 109658 590698 109894
rect 590142 109338 590378 109574
rect 590462 109338 590698 109574
rect 590142 69658 590378 69894
rect 590462 69658 590698 69894
rect 590142 69338 590378 69574
rect 590462 69338 590698 69574
rect 590142 29658 590378 29894
rect 590462 29658 590698 29894
rect 590142 29338 590378 29574
rect 590462 29338 590698 29574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 693378 591338 693614
rect 591422 693378 591658 693614
rect 591102 693058 591338 693294
rect 591422 693058 591658 693294
rect 591102 653378 591338 653614
rect 591422 653378 591658 653614
rect 591102 653058 591338 653294
rect 591422 653058 591658 653294
rect 591102 613378 591338 613614
rect 591422 613378 591658 613614
rect 591102 613058 591338 613294
rect 591422 613058 591658 613294
rect 591102 573378 591338 573614
rect 591422 573378 591658 573614
rect 591102 573058 591338 573294
rect 591422 573058 591658 573294
rect 591102 533378 591338 533614
rect 591422 533378 591658 533614
rect 591102 533058 591338 533294
rect 591422 533058 591658 533294
rect 591102 493378 591338 493614
rect 591422 493378 591658 493614
rect 591102 493058 591338 493294
rect 591422 493058 591658 493294
rect 591102 453378 591338 453614
rect 591422 453378 591658 453614
rect 591102 453058 591338 453294
rect 591422 453058 591658 453294
rect 591102 413378 591338 413614
rect 591422 413378 591658 413614
rect 591102 413058 591338 413294
rect 591422 413058 591658 413294
rect 591102 373378 591338 373614
rect 591422 373378 591658 373614
rect 591102 373058 591338 373294
rect 591422 373058 591658 373294
rect 591102 333378 591338 333614
rect 591422 333378 591658 333614
rect 591102 333058 591338 333294
rect 591422 333058 591658 333294
rect 591102 293378 591338 293614
rect 591422 293378 591658 293614
rect 591102 293058 591338 293294
rect 591422 293058 591658 293294
rect 591102 253378 591338 253614
rect 591422 253378 591658 253614
rect 591102 253058 591338 253294
rect 591422 253058 591658 253294
rect 591102 213378 591338 213614
rect 591422 213378 591658 213614
rect 591102 213058 591338 213294
rect 591422 213058 591658 213294
rect 591102 173378 591338 173614
rect 591422 173378 591658 173614
rect 591102 173058 591338 173294
rect 591422 173058 591658 173294
rect 591102 133378 591338 133614
rect 591422 133378 591658 133614
rect 591102 133058 591338 133294
rect 591422 133058 591658 133294
rect 591102 93378 591338 93614
rect 591422 93378 591658 93614
rect 591102 93058 591338 93294
rect 591422 93058 591658 93294
rect 591102 53378 591338 53614
rect 591422 53378 591658 53614
rect 591102 53058 591338 53294
rect 591422 53058 591658 53294
rect 591102 13378 591338 13614
rect 591422 13378 591658 13614
rect 591102 13058 591338 13294
rect 591422 13058 591658 13294
rect 571986 -6342 572222 -6106
rect 572306 -6342 572542 -6106
rect 571986 -6662 572222 -6426
rect 572306 -6662 572542 -6426
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 673378 592298 673614
rect 592382 673378 592618 673614
rect 592062 673058 592298 673294
rect 592382 673058 592618 673294
rect 592062 633378 592298 633614
rect 592382 633378 592618 633614
rect 592062 633058 592298 633294
rect 592382 633058 592618 633294
rect 592062 593378 592298 593614
rect 592382 593378 592618 593614
rect 592062 593058 592298 593294
rect 592382 593058 592618 593294
rect 592062 553378 592298 553614
rect 592382 553378 592618 553614
rect 592062 553058 592298 553294
rect 592382 553058 592618 553294
rect 592062 513378 592298 513614
rect 592382 513378 592618 513614
rect 592062 513058 592298 513294
rect 592382 513058 592618 513294
rect 592062 473378 592298 473614
rect 592382 473378 592618 473614
rect 592062 473058 592298 473294
rect 592382 473058 592618 473294
rect 592062 433378 592298 433614
rect 592382 433378 592618 433614
rect 592062 433058 592298 433294
rect 592382 433058 592618 433294
rect 592062 393378 592298 393614
rect 592382 393378 592618 393614
rect 592062 393058 592298 393294
rect 592382 393058 592618 393294
rect 592062 353378 592298 353614
rect 592382 353378 592618 353614
rect 592062 353058 592298 353294
rect 592382 353058 592618 353294
rect 592062 313378 592298 313614
rect 592382 313378 592618 313614
rect 592062 313058 592298 313294
rect 592382 313058 592618 313294
rect 592062 273378 592298 273614
rect 592382 273378 592618 273614
rect 592062 273058 592298 273294
rect 592382 273058 592618 273294
rect 592062 233378 592298 233614
rect 592382 233378 592618 233614
rect 592062 233058 592298 233294
rect 592382 233058 592618 233294
rect 592062 193378 592298 193614
rect 592382 193378 592618 193614
rect 592062 193058 592298 193294
rect 592382 193058 592618 193294
rect 592062 153378 592298 153614
rect 592382 153378 592618 153614
rect 592062 153058 592298 153294
rect 592382 153058 592618 153294
rect 592062 113378 592298 113614
rect 592382 113378 592618 113614
rect 592062 113058 592298 113294
rect 592382 113058 592618 113294
rect 592062 73378 592298 73614
rect 592382 73378 592618 73614
rect 592062 73058 592298 73294
rect 592382 73058 592618 73294
rect 592062 33378 592298 33614
rect 592382 33378 592618 33614
rect 592062 33058 592298 33294
rect 592382 33058 592618 33294
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 31986 711558
rect 32222 711322 32306 711558
rect 32542 711322 71986 711558
rect 72222 711322 72306 711558
rect 72542 711322 111986 711558
rect 112222 711322 112306 711558
rect 112542 711322 151986 711558
rect 152222 711322 152306 711558
rect 152542 711322 191986 711558
rect 192222 711322 192306 711558
rect 192542 711322 231986 711558
rect 232222 711322 232306 711558
rect 232542 711322 271986 711558
rect 272222 711322 272306 711558
rect 272542 711322 311986 711558
rect 312222 711322 312306 711558
rect 312542 711322 351986 711558
rect 352222 711322 352306 711558
rect 352542 711322 391986 711558
rect 392222 711322 392306 711558
rect 392542 711322 431986 711558
rect 432222 711322 432306 711558
rect 432542 711322 471986 711558
rect 472222 711322 472306 711558
rect 472542 711322 511986 711558
rect 512222 711322 512306 711558
rect 512542 711322 551986 711558
rect 552222 711322 552306 711558
rect 552542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 31986 711238
rect 32222 711002 32306 711238
rect 32542 711002 71986 711238
rect 72222 711002 72306 711238
rect 72542 711002 111986 711238
rect 112222 711002 112306 711238
rect 112542 711002 151986 711238
rect 152222 711002 152306 711238
rect 152542 711002 191986 711238
rect 192222 711002 192306 711238
rect 192542 711002 231986 711238
rect 232222 711002 232306 711238
rect 232542 711002 271986 711238
rect 272222 711002 272306 711238
rect 272542 711002 311986 711238
rect 312222 711002 312306 711238
rect 312542 711002 351986 711238
rect 352222 711002 352306 711238
rect 352542 711002 391986 711238
rect 392222 711002 392306 711238
rect 392542 711002 431986 711238
rect 432222 711002 432306 711238
rect 432542 711002 471986 711238
rect 472222 711002 472306 711238
rect 472542 711002 511986 711238
rect 512222 711002 512306 711238
rect 512542 711002 551986 711238
rect 552222 711002 552306 711238
rect 552542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 11986 710598
rect 12222 710362 12306 710598
rect 12542 710362 51986 710598
rect 52222 710362 52306 710598
rect 52542 710362 91986 710598
rect 92222 710362 92306 710598
rect 92542 710362 131986 710598
rect 132222 710362 132306 710598
rect 132542 710362 171986 710598
rect 172222 710362 172306 710598
rect 172542 710362 211986 710598
rect 212222 710362 212306 710598
rect 212542 710362 251986 710598
rect 252222 710362 252306 710598
rect 252542 710362 291986 710598
rect 292222 710362 292306 710598
rect 292542 710362 331986 710598
rect 332222 710362 332306 710598
rect 332542 710362 371986 710598
rect 372222 710362 372306 710598
rect 372542 710362 411986 710598
rect 412222 710362 412306 710598
rect 412542 710362 451986 710598
rect 452222 710362 452306 710598
rect 452542 710362 491986 710598
rect 492222 710362 492306 710598
rect 492542 710362 531986 710598
rect 532222 710362 532306 710598
rect 532542 710362 571986 710598
rect 572222 710362 572306 710598
rect 572542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 11986 710278
rect 12222 710042 12306 710278
rect 12542 710042 51986 710278
rect 52222 710042 52306 710278
rect 52542 710042 91986 710278
rect 92222 710042 92306 710278
rect 92542 710042 131986 710278
rect 132222 710042 132306 710278
rect 132542 710042 171986 710278
rect 172222 710042 172306 710278
rect 172542 710042 211986 710278
rect 212222 710042 212306 710278
rect 212542 710042 251986 710278
rect 252222 710042 252306 710278
rect 252542 710042 291986 710278
rect 292222 710042 292306 710278
rect 292542 710042 331986 710278
rect 332222 710042 332306 710278
rect 332542 710042 371986 710278
rect 372222 710042 372306 710278
rect 372542 710042 411986 710278
rect 412222 710042 412306 710278
rect 412542 710042 451986 710278
rect 452222 710042 452306 710278
rect 452542 710042 491986 710278
rect 492222 710042 492306 710278
rect 492542 710042 531986 710278
rect 532222 710042 532306 710278
rect 532542 710042 571986 710278
rect 572222 710042 572306 710278
rect 572542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 28266 709638
rect 28502 709402 28586 709638
rect 28822 709402 68266 709638
rect 68502 709402 68586 709638
rect 68822 709402 108266 709638
rect 108502 709402 108586 709638
rect 108822 709402 148266 709638
rect 148502 709402 148586 709638
rect 148822 709402 188266 709638
rect 188502 709402 188586 709638
rect 188822 709402 228266 709638
rect 228502 709402 228586 709638
rect 228822 709402 268266 709638
rect 268502 709402 268586 709638
rect 268822 709402 308266 709638
rect 308502 709402 308586 709638
rect 308822 709402 348266 709638
rect 348502 709402 348586 709638
rect 348822 709402 388266 709638
rect 388502 709402 388586 709638
rect 388822 709402 428266 709638
rect 428502 709402 428586 709638
rect 428822 709402 468266 709638
rect 468502 709402 468586 709638
rect 468822 709402 508266 709638
rect 508502 709402 508586 709638
rect 508822 709402 548266 709638
rect 548502 709402 548586 709638
rect 548822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 28266 709318
rect 28502 709082 28586 709318
rect 28822 709082 68266 709318
rect 68502 709082 68586 709318
rect 68822 709082 108266 709318
rect 108502 709082 108586 709318
rect 108822 709082 148266 709318
rect 148502 709082 148586 709318
rect 148822 709082 188266 709318
rect 188502 709082 188586 709318
rect 188822 709082 228266 709318
rect 228502 709082 228586 709318
rect 228822 709082 268266 709318
rect 268502 709082 268586 709318
rect 268822 709082 308266 709318
rect 308502 709082 308586 709318
rect 308822 709082 348266 709318
rect 348502 709082 348586 709318
rect 348822 709082 388266 709318
rect 388502 709082 388586 709318
rect 388822 709082 428266 709318
rect 428502 709082 428586 709318
rect 428822 709082 468266 709318
rect 468502 709082 468586 709318
rect 468822 709082 508266 709318
rect 508502 709082 508586 709318
rect 508822 709082 548266 709318
rect 548502 709082 548586 709318
rect 548822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 8266 708678
rect 8502 708442 8586 708678
rect 8822 708442 48266 708678
rect 48502 708442 48586 708678
rect 48822 708442 88266 708678
rect 88502 708442 88586 708678
rect 88822 708442 128266 708678
rect 128502 708442 128586 708678
rect 128822 708442 168266 708678
rect 168502 708442 168586 708678
rect 168822 708442 208266 708678
rect 208502 708442 208586 708678
rect 208822 708442 248266 708678
rect 248502 708442 248586 708678
rect 248822 708442 288266 708678
rect 288502 708442 288586 708678
rect 288822 708442 328266 708678
rect 328502 708442 328586 708678
rect 328822 708442 368266 708678
rect 368502 708442 368586 708678
rect 368822 708442 408266 708678
rect 408502 708442 408586 708678
rect 408822 708442 448266 708678
rect 448502 708442 448586 708678
rect 448822 708442 488266 708678
rect 488502 708442 488586 708678
rect 488822 708442 528266 708678
rect 528502 708442 528586 708678
rect 528822 708442 568266 708678
rect 568502 708442 568586 708678
rect 568822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 8266 708358
rect 8502 708122 8586 708358
rect 8822 708122 48266 708358
rect 48502 708122 48586 708358
rect 48822 708122 88266 708358
rect 88502 708122 88586 708358
rect 88822 708122 128266 708358
rect 128502 708122 128586 708358
rect 128822 708122 168266 708358
rect 168502 708122 168586 708358
rect 168822 708122 208266 708358
rect 208502 708122 208586 708358
rect 208822 708122 248266 708358
rect 248502 708122 248586 708358
rect 248822 708122 288266 708358
rect 288502 708122 288586 708358
rect 288822 708122 328266 708358
rect 328502 708122 328586 708358
rect 328822 708122 368266 708358
rect 368502 708122 368586 708358
rect 368822 708122 408266 708358
rect 408502 708122 408586 708358
rect 408822 708122 448266 708358
rect 448502 708122 448586 708358
rect 448822 708122 488266 708358
rect 488502 708122 488586 708358
rect 488822 708122 528266 708358
rect 528502 708122 528586 708358
rect 528822 708122 568266 708358
rect 568502 708122 568586 708358
rect 568822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 24546 707718
rect 24782 707482 24866 707718
rect 25102 707482 64546 707718
rect 64782 707482 64866 707718
rect 65102 707482 104546 707718
rect 104782 707482 104866 707718
rect 105102 707482 144546 707718
rect 144782 707482 144866 707718
rect 145102 707482 184546 707718
rect 184782 707482 184866 707718
rect 185102 707482 224546 707718
rect 224782 707482 224866 707718
rect 225102 707482 264546 707718
rect 264782 707482 264866 707718
rect 265102 707482 304546 707718
rect 304782 707482 304866 707718
rect 305102 707482 344546 707718
rect 344782 707482 344866 707718
rect 345102 707482 384546 707718
rect 384782 707482 384866 707718
rect 385102 707482 424546 707718
rect 424782 707482 424866 707718
rect 425102 707482 464546 707718
rect 464782 707482 464866 707718
rect 465102 707482 504546 707718
rect 504782 707482 504866 707718
rect 505102 707482 544546 707718
rect 544782 707482 544866 707718
rect 545102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 24546 707398
rect 24782 707162 24866 707398
rect 25102 707162 64546 707398
rect 64782 707162 64866 707398
rect 65102 707162 104546 707398
rect 104782 707162 104866 707398
rect 105102 707162 144546 707398
rect 144782 707162 144866 707398
rect 145102 707162 184546 707398
rect 184782 707162 184866 707398
rect 185102 707162 224546 707398
rect 224782 707162 224866 707398
rect 225102 707162 264546 707398
rect 264782 707162 264866 707398
rect 265102 707162 304546 707398
rect 304782 707162 304866 707398
rect 305102 707162 344546 707398
rect 344782 707162 344866 707398
rect 345102 707162 384546 707398
rect 384782 707162 384866 707398
rect 385102 707162 424546 707398
rect 424782 707162 424866 707398
rect 425102 707162 464546 707398
rect 464782 707162 464866 707398
rect 465102 707162 504546 707398
rect 504782 707162 504866 707398
rect 505102 707162 544546 707398
rect 544782 707162 544866 707398
rect 545102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 4546 706758
rect 4782 706522 4866 706758
rect 5102 706522 44546 706758
rect 44782 706522 44866 706758
rect 45102 706522 84546 706758
rect 84782 706522 84866 706758
rect 85102 706522 124546 706758
rect 124782 706522 124866 706758
rect 125102 706522 164546 706758
rect 164782 706522 164866 706758
rect 165102 706522 204546 706758
rect 204782 706522 204866 706758
rect 205102 706522 244546 706758
rect 244782 706522 244866 706758
rect 245102 706522 284546 706758
rect 284782 706522 284866 706758
rect 285102 706522 324546 706758
rect 324782 706522 324866 706758
rect 325102 706522 364546 706758
rect 364782 706522 364866 706758
rect 365102 706522 404546 706758
rect 404782 706522 404866 706758
rect 405102 706522 444546 706758
rect 444782 706522 444866 706758
rect 445102 706522 484546 706758
rect 484782 706522 484866 706758
rect 485102 706522 524546 706758
rect 524782 706522 524866 706758
rect 525102 706522 564546 706758
rect 564782 706522 564866 706758
rect 565102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 4546 706438
rect 4782 706202 4866 706438
rect 5102 706202 44546 706438
rect 44782 706202 44866 706438
rect 45102 706202 84546 706438
rect 84782 706202 84866 706438
rect 85102 706202 124546 706438
rect 124782 706202 124866 706438
rect 125102 706202 164546 706438
rect 164782 706202 164866 706438
rect 165102 706202 204546 706438
rect 204782 706202 204866 706438
rect 205102 706202 244546 706438
rect 244782 706202 244866 706438
rect 245102 706202 284546 706438
rect 284782 706202 284866 706438
rect 285102 706202 324546 706438
rect 324782 706202 324866 706438
rect 325102 706202 364546 706438
rect 364782 706202 364866 706438
rect 365102 706202 404546 706438
rect 404782 706202 404866 706438
rect 405102 706202 444546 706438
rect 444782 706202 444866 706438
rect 445102 706202 484546 706438
rect 484782 706202 484866 706438
rect 485102 706202 524546 706438
rect 524782 706202 524866 706438
rect 525102 706202 564546 706438
rect 564782 706202 564866 706438
rect 565102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 20826 705798
rect 21062 705562 21146 705798
rect 21382 705562 60826 705798
rect 61062 705562 61146 705798
rect 61382 705562 100826 705798
rect 101062 705562 101146 705798
rect 101382 705562 140826 705798
rect 141062 705562 141146 705798
rect 141382 705562 180826 705798
rect 181062 705562 181146 705798
rect 181382 705562 220826 705798
rect 221062 705562 221146 705798
rect 221382 705562 260826 705798
rect 261062 705562 261146 705798
rect 261382 705562 300826 705798
rect 301062 705562 301146 705798
rect 301382 705562 340826 705798
rect 341062 705562 341146 705798
rect 341382 705562 380826 705798
rect 381062 705562 381146 705798
rect 381382 705562 420826 705798
rect 421062 705562 421146 705798
rect 421382 705562 460826 705798
rect 461062 705562 461146 705798
rect 461382 705562 500826 705798
rect 501062 705562 501146 705798
rect 501382 705562 540826 705798
rect 541062 705562 541146 705798
rect 541382 705562 580826 705798
rect 581062 705562 581146 705798
rect 581382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 20826 705478
rect 21062 705242 21146 705478
rect 21382 705242 60826 705478
rect 61062 705242 61146 705478
rect 61382 705242 100826 705478
rect 101062 705242 101146 705478
rect 101382 705242 140826 705478
rect 141062 705242 141146 705478
rect 141382 705242 180826 705478
rect 181062 705242 181146 705478
rect 181382 705242 220826 705478
rect 221062 705242 221146 705478
rect 221382 705242 260826 705478
rect 261062 705242 261146 705478
rect 261382 705242 300826 705478
rect 301062 705242 301146 705478
rect 301382 705242 340826 705478
rect 341062 705242 341146 705478
rect 341382 705242 380826 705478
rect 381062 705242 381146 705478
rect 381382 705242 420826 705478
rect 421062 705242 421146 705478
rect 421382 705242 460826 705478
rect 461062 705242 461146 705478
rect 461382 705242 500826 705478
rect 501062 705242 501146 705478
rect 501382 705242 540826 705478
rect 541062 705242 541146 705478
rect 541382 705242 580826 705478
rect 581062 705242 581146 705478
rect 581382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 826 704838
rect 1062 704602 1146 704838
rect 1382 704602 40826 704838
rect 41062 704602 41146 704838
rect 41382 704602 80826 704838
rect 81062 704602 81146 704838
rect 81382 704602 120826 704838
rect 121062 704602 121146 704838
rect 121382 704602 160826 704838
rect 161062 704602 161146 704838
rect 161382 704602 200826 704838
rect 201062 704602 201146 704838
rect 201382 704602 240826 704838
rect 241062 704602 241146 704838
rect 241382 704602 280826 704838
rect 281062 704602 281146 704838
rect 281382 704602 320826 704838
rect 321062 704602 321146 704838
rect 321382 704602 360826 704838
rect 361062 704602 361146 704838
rect 361382 704602 400826 704838
rect 401062 704602 401146 704838
rect 401382 704602 440826 704838
rect 441062 704602 441146 704838
rect 441382 704602 480826 704838
rect 481062 704602 481146 704838
rect 481382 704602 520826 704838
rect 521062 704602 521146 704838
rect 521382 704602 560826 704838
rect 561062 704602 561146 704838
rect 561382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 826 704518
rect 1062 704282 1146 704518
rect 1382 704282 40826 704518
rect 41062 704282 41146 704518
rect 41382 704282 80826 704518
rect 81062 704282 81146 704518
rect 81382 704282 120826 704518
rect 121062 704282 121146 704518
rect 121382 704282 160826 704518
rect 161062 704282 161146 704518
rect 161382 704282 200826 704518
rect 201062 704282 201146 704518
rect 201382 704282 240826 704518
rect 241062 704282 241146 704518
rect 241382 704282 280826 704518
rect 281062 704282 281146 704518
rect 281382 704282 320826 704518
rect 321062 704282 321146 704518
rect 321382 704282 360826 704518
rect 361062 704282 361146 704518
rect 361382 704282 400826 704518
rect 401062 704282 401146 704518
rect 401382 704282 440826 704518
rect 441062 704282 441146 704518
rect 441382 704282 480826 704518
rect 481062 704282 481146 704518
rect 481382 704282 520826 704518
rect 521062 704282 521146 704518
rect 521382 704282 560826 704518
rect 561062 704282 561146 704518
rect 561382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 693614 592650 693646
rect -8726 693378 -7734 693614
rect -7498 693378 -7414 693614
rect -7178 693378 11986 693614
rect 12222 693378 12306 693614
rect 12542 693378 51986 693614
rect 52222 693378 52306 693614
rect 52542 693378 91986 693614
rect 92222 693378 92306 693614
rect 92542 693378 131986 693614
rect 132222 693378 132306 693614
rect 132542 693378 171986 693614
rect 172222 693378 172306 693614
rect 172542 693378 211986 693614
rect 212222 693378 212306 693614
rect 212542 693378 251986 693614
rect 252222 693378 252306 693614
rect 252542 693378 291986 693614
rect 292222 693378 292306 693614
rect 292542 693378 331986 693614
rect 332222 693378 332306 693614
rect 332542 693378 371986 693614
rect 372222 693378 372306 693614
rect 372542 693378 411986 693614
rect 412222 693378 412306 693614
rect 412542 693378 451986 693614
rect 452222 693378 452306 693614
rect 452542 693378 491986 693614
rect 492222 693378 492306 693614
rect 492542 693378 531986 693614
rect 532222 693378 532306 693614
rect 532542 693378 571986 693614
rect 572222 693378 572306 693614
rect 572542 693378 591102 693614
rect 591338 693378 591422 693614
rect 591658 693378 592650 693614
rect -8726 693294 592650 693378
rect -8726 693058 -7734 693294
rect -7498 693058 -7414 693294
rect -7178 693058 11986 693294
rect 12222 693058 12306 693294
rect 12542 693058 51986 693294
rect 52222 693058 52306 693294
rect 52542 693058 91986 693294
rect 92222 693058 92306 693294
rect 92542 693058 131986 693294
rect 132222 693058 132306 693294
rect 132542 693058 171986 693294
rect 172222 693058 172306 693294
rect 172542 693058 211986 693294
rect 212222 693058 212306 693294
rect 212542 693058 251986 693294
rect 252222 693058 252306 693294
rect 252542 693058 291986 693294
rect 292222 693058 292306 693294
rect 292542 693058 331986 693294
rect 332222 693058 332306 693294
rect 332542 693058 371986 693294
rect 372222 693058 372306 693294
rect 372542 693058 411986 693294
rect 412222 693058 412306 693294
rect 412542 693058 451986 693294
rect 452222 693058 452306 693294
rect 452542 693058 491986 693294
rect 492222 693058 492306 693294
rect 492542 693058 531986 693294
rect 532222 693058 532306 693294
rect 532542 693058 571986 693294
rect 572222 693058 572306 693294
rect 572542 693058 591102 693294
rect 591338 693058 591422 693294
rect 591658 693058 592650 693294
rect -8726 693026 592650 693058
rect -6806 689894 590730 689926
rect -6806 689658 -5814 689894
rect -5578 689658 -5494 689894
rect -5258 689658 8266 689894
rect 8502 689658 8586 689894
rect 8822 689658 48266 689894
rect 48502 689658 48586 689894
rect 48822 689658 88266 689894
rect 88502 689658 88586 689894
rect 88822 689658 128266 689894
rect 128502 689658 128586 689894
rect 128822 689658 168266 689894
rect 168502 689658 168586 689894
rect 168822 689658 208266 689894
rect 208502 689658 208586 689894
rect 208822 689658 248266 689894
rect 248502 689658 248586 689894
rect 248822 689658 288266 689894
rect 288502 689658 288586 689894
rect 288822 689658 328266 689894
rect 328502 689658 328586 689894
rect 328822 689658 368266 689894
rect 368502 689658 368586 689894
rect 368822 689658 408266 689894
rect 408502 689658 408586 689894
rect 408822 689658 448266 689894
rect 448502 689658 448586 689894
rect 448822 689658 488266 689894
rect 488502 689658 488586 689894
rect 488822 689658 528266 689894
rect 528502 689658 528586 689894
rect 528822 689658 568266 689894
rect 568502 689658 568586 689894
rect 568822 689658 589182 689894
rect 589418 689658 589502 689894
rect 589738 689658 590730 689894
rect -6806 689574 590730 689658
rect -6806 689338 -5814 689574
rect -5578 689338 -5494 689574
rect -5258 689338 8266 689574
rect 8502 689338 8586 689574
rect 8822 689338 48266 689574
rect 48502 689338 48586 689574
rect 48822 689338 88266 689574
rect 88502 689338 88586 689574
rect 88822 689338 128266 689574
rect 128502 689338 128586 689574
rect 128822 689338 168266 689574
rect 168502 689338 168586 689574
rect 168822 689338 208266 689574
rect 208502 689338 208586 689574
rect 208822 689338 248266 689574
rect 248502 689338 248586 689574
rect 248822 689338 288266 689574
rect 288502 689338 288586 689574
rect 288822 689338 328266 689574
rect 328502 689338 328586 689574
rect 328822 689338 368266 689574
rect 368502 689338 368586 689574
rect 368822 689338 408266 689574
rect 408502 689338 408586 689574
rect 408822 689338 448266 689574
rect 448502 689338 448586 689574
rect 448822 689338 488266 689574
rect 488502 689338 488586 689574
rect 488822 689338 528266 689574
rect 528502 689338 528586 689574
rect 528822 689338 568266 689574
rect 568502 689338 568586 689574
rect 568822 689338 589182 689574
rect 589418 689338 589502 689574
rect 589738 689338 590730 689574
rect -6806 689306 590730 689338
rect -4886 686174 588810 686206
rect -4886 685938 -3894 686174
rect -3658 685938 -3574 686174
rect -3338 685938 4546 686174
rect 4782 685938 4866 686174
rect 5102 685938 44546 686174
rect 44782 685938 44866 686174
rect 45102 685938 84546 686174
rect 84782 685938 84866 686174
rect 85102 685938 124546 686174
rect 124782 685938 124866 686174
rect 125102 685938 164546 686174
rect 164782 685938 164866 686174
rect 165102 685938 204546 686174
rect 204782 685938 204866 686174
rect 205102 685938 244546 686174
rect 244782 685938 244866 686174
rect 245102 685938 284546 686174
rect 284782 685938 284866 686174
rect 285102 685938 324546 686174
rect 324782 685938 324866 686174
rect 325102 685938 364546 686174
rect 364782 685938 364866 686174
rect 365102 685938 404546 686174
rect 404782 685938 404866 686174
rect 405102 685938 444546 686174
rect 444782 685938 444866 686174
rect 445102 685938 484546 686174
rect 484782 685938 484866 686174
rect 485102 685938 524546 686174
rect 524782 685938 524866 686174
rect 525102 685938 564546 686174
rect 564782 685938 564866 686174
rect 565102 685938 587262 686174
rect 587498 685938 587582 686174
rect 587818 685938 588810 686174
rect -4886 685854 588810 685938
rect -4886 685618 -3894 685854
rect -3658 685618 -3574 685854
rect -3338 685618 4546 685854
rect 4782 685618 4866 685854
rect 5102 685618 44546 685854
rect 44782 685618 44866 685854
rect 45102 685618 84546 685854
rect 84782 685618 84866 685854
rect 85102 685618 124546 685854
rect 124782 685618 124866 685854
rect 125102 685618 164546 685854
rect 164782 685618 164866 685854
rect 165102 685618 204546 685854
rect 204782 685618 204866 685854
rect 205102 685618 244546 685854
rect 244782 685618 244866 685854
rect 245102 685618 284546 685854
rect 284782 685618 284866 685854
rect 285102 685618 324546 685854
rect 324782 685618 324866 685854
rect 325102 685618 364546 685854
rect 364782 685618 364866 685854
rect 365102 685618 404546 685854
rect 404782 685618 404866 685854
rect 405102 685618 444546 685854
rect 444782 685618 444866 685854
rect 445102 685618 484546 685854
rect 484782 685618 484866 685854
rect 485102 685618 524546 685854
rect 524782 685618 524866 685854
rect 525102 685618 564546 685854
rect 564782 685618 564866 685854
rect 565102 685618 587262 685854
rect 587498 685618 587582 685854
rect 587818 685618 588810 685854
rect -4886 685586 588810 685618
rect -2966 682454 586890 682486
rect -2966 682218 -1974 682454
rect -1738 682218 -1654 682454
rect -1418 682218 826 682454
rect 1062 682218 1146 682454
rect 1382 682218 40826 682454
rect 41062 682218 41146 682454
rect 41382 682218 80826 682454
rect 81062 682218 81146 682454
rect 81382 682218 120826 682454
rect 121062 682218 121146 682454
rect 121382 682218 160826 682454
rect 161062 682218 161146 682454
rect 161382 682218 200826 682454
rect 201062 682218 201146 682454
rect 201382 682218 240826 682454
rect 241062 682218 241146 682454
rect 241382 682218 280826 682454
rect 281062 682218 281146 682454
rect 281382 682218 320826 682454
rect 321062 682218 321146 682454
rect 321382 682218 360826 682454
rect 361062 682218 361146 682454
rect 361382 682218 400826 682454
rect 401062 682218 401146 682454
rect 401382 682218 440826 682454
rect 441062 682218 441146 682454
rect 441382 682218 480826 682454
rect 481062 682218 481146 682454
rect 481382 682218 520826 682454
rect 521062 682218 521146 682454
rect 521382 682218 560826 682454
rect 561062 682218 561146 682454
rect 561382 682218 585342 682454
rect 585578 682218 585662 682454
rect 585898 682218 586890 682454
rect -2966 682134 586890 682218
rect -2966 681898 -1974 682134
rect -1738 681898 -1654 682134
rect -1418 681898 826 682134
rect 1062 681898 1146 682134
rect 1382 681898 40826 682134
rect 41062 681898 41146 682134
rect 41382 681898 80826 682134
rect 81062 681898 81146 682134
rect 81382 681898 120826 682134
rect 121062 681898 121146 682134
rect 121382 681898 160826 682134
rect 161062 681898 161146 682134
rect 161382 681898 200826 682134
rect 201062 681898 201146 682134
rect 201382 681898 240826 682134
rect 241062 681898 241146 682134
rect 241382 681898 280826 682134
rect 281062 681898 281146 682134
rect 281382 681898 320826 682134
rect 321062 681898 321146 682134
rect 321382 681898 360826 682134
rect 361062 681898 361146 682134
rect 361382 681898 400826 682134
rect 401062 681898 401146 682134
rect 401382 681898 440826 682134
rect 441062 681898 441146 682134
rect 441382 681898 480826 682134
rect 481062 681898 481146 682134
rect 481382 681898 520826 682134
rect 521062 681898 521146 682134
rect 521382 681898 560826 682134
rect 561062 681898 561146 682134
rect 561382 681898 585342 682134
rect 585578 681898 585662 682134
rect 585898 681898 586890 682134
rect -2966 681866 586890 681898
rect -8726 673614 592650 673646
rect -8726 673378 -8694 673614
rect -8458 673378 -8374 673614
rect -8138 673378 31986 673614
rect 32222 673378 32306 673614
rect 32542 673378 71986 673614
rect 72222 673378 72306 673614
rect 72542 673378 111986 673614
rect 112222 673378 112306 673614
rect 112542 673378 151986 673614
rect 152222 673378 152306 673614
rect 152542 673378 191986 673614
rect 192222 673378 192306 673614
rect 192542 673378 231986 673614
rect 232222 673378 232306 673614
rect 232542 673378 271986 673614
rect 272222 673378 272306 673614
rect 272542 673378 311986 673614
rect 312222 673378 312306 673614
rect 312542 673378 351986 673614
rect 352222 673378 352306 673614
rect 352542 673378 391986 673614
rect 392222 673378 392306 673614
rect 392542 673378 431986 673614
rect 432222 673378 432306 673614
rect 432542 673378 471986 673614
rect 472222 673378 472306 673614
rect 472542 673378 511986 673614
rect 512222 673378 512306 673614
rect 512542 673378 551986 673614
rect 552222 673378 552306 673614
rect 552542 673378 592062 673614
rect 592298 673378 592382 673614
rect 592618 673378 592650 673614
rect -8726 673294 592650 673378
rect -8726 673058 -8694 673294
rect -8458 673058 -8374 673294
rect -8138 673058 31986 673294
rect 32222 673058 32306 673294
rect 32542 673058 71986 673294
rect 72222 673058 72306 673294
rect 72542 673058 111986 673294
rect 112222 673058 112306 673294
rect 112542 673058 151986 673294
rect 152222 673058 152306 673294
rect 152542 673058 191986 673294
rect 192222 673058 192306 673294
rect 192542 673058 231986 673294
rect 232222 673058 232306 673294
rect 232542 673058 271986 673294
rect 272222 673058 272306 673294
rect 272542 673058 311986 673294
rect 312222 673058 312306 673294
rect 312542 673058 351986 673294
rect 352222 673058 352306 673294
rect 352542 673058 391986 673294
rect 392222 673058 392306 673294
rect 392542 673058 431986 673294
rect 432222 673058 432306 673294
rect 432542 673058 471986 673294
rect 472222 673058 472306 673294
rect 472542 673058 511986 673294
rect 512222 673058 512306 673294
rect 512542 673058 551986 673294
rect 552222 673058 552306 673294
rect 552542 673058 592062 673294
rect 592298 673058 592382 673294
rect 592618 673058 592650 673294
rect -8726 673026 592650 673058
rect -6806 669894 590730 669926
rect -6806 669658 -6774 669894
rect -6538 669658 -6454 669894
rect -6218 669658 28266 669894
rect 28502 669658 28586 669894
rect 28822 669658 68266 669894
rect 68502 669658 68586 669894
rect 68822 669658 108266 669894
rect 108502 669658 108586 669894
rect 108822 669658 148266 669894
rect 148502 669658 148586 669894
rect 148822 669658 188266 669894
rect 188502 669658 188586 669894
rect 188822 669658 228266 669894
rect 228502 669658 228586 669894
rect 228822 669658 268266 669894
rect 268502 669658 268586 669894
rect 268822 669658 308266 669894
rect 308502 669658 308586 669894
rect 308822 669658 348266 669894
rect 348502 669658 348586 669894
rect 348822 669658 388266 669894
rect 388502 669658 388586 669894
rect 388822 669658 428266 669894
rect 428502 669658 428586 669894
rect 428822 669658 468266 669894
rect 468502 669658 468586 669894
rect 468822 669658 508266 669894
rect 508502 669658 508586 669894
rect 508822 669658 548266 669894
rect 548502 669658 548586 669894
rect 548822 669658 590142 669894
rect 590378 669658 590462 669894
rect 590698 669658 590730 669894
rect -6806 669574 590730 669658
rect -6806 669338 -6774 669574
rect -6538 669338 -6454 669574
rect -6218 669338 28266 669574
rect 28502 669338 28586 669574
rect 28822 669338 68266 669574
rect 68502 669338 68586 669574
rect 68822 669338 108266 669574
rect 108502 669338 108586 669574
rect 108822 669338 148266 669574
rect 148502 669338 148586 669574
rect 148822 669338 188266 669574
rect 188502 669338 188586 669574
rect 188822 669338 228266 669574
rect 228502 669338 228586 669574
rect 228822 669338 268266 669574
rect 268502 669338 268586 669574
rect 268822 669338 308266 669574
rect 308502 669338 308586 669574
rect 308822 669338 348266 669574
rect 348502 669338 348586 669574
rect 348822 669338 388266 669574
rect 388502 669338 388586 669574
rect 388822 669338 428266 669574
rect 428502 669338 428586 669574
rect 428822 669338 468266 669574
rect 468502 669338 468586 669574
rect 468822 669338 508266 669574
rect 508502 669338 508586 669574
rect 508822 669338 548266 669574
rect 548502 669338 548586 669574
rect 548822 669338 590142 669574
rect 590378 669338 590462 669574
rect 590698 669338 590730 669574
rect -6806 669306 590730 669338
rect -4886 666174 588810 666206
rect -4886 665938 -4854 666174
rect -4618 665938 -4534 666174
rect -4298 665938 24546 666174
rect 24782 665938 24866 666174
rect 25102 665938 64546 666174
rect 64782 665938 64866 666174
rect 65102 665938 104546 666174
rect 104782 665938 104866 666174
rect 105102 665938 144546 666174
rect 144782 665938 144866 666174
rect 145102 665938 184546 666174
rect 184782 665938 184866 666174
rect 185102 665938 224546 666174
rect 224782 665938 224866 666174
rect 225102 665938 264546 666174
rect 264782 665938 264866 666174
rect 265102 665938 304546 666174
rect 304782 665938 304866 666174
rect 305102 665938 344546 666174
rect 344782 665938 344866 666174
rect 345102 665938 384546 666174
rect 384782 665938 384866 666174
rect 385102 665938 424546 666174
rect 424782 665938 424866 666174
rect 425102 665938 464546 666174
rect 464782 665938 464866 666174
rect 465102 665938 504546 666174
rect 504782 665938 504866 666174
rect 505102 665938 544546 666174
rect 544782 665938 544866 666174
rect 545102 665938 588222 666174
rect 588458 665938 588542 666174
rect 588778 665938 588810 666174
rect -4886 665854 588810 665938
rect -4886 665618 -4854 665854
rect -4618 665618 -4534 665854
rect -4298 665618 24546 665854
rect 24782 665618 24866 665854
rect 25102 665618 64546 665854
rect 64782 665618 64866 665854
rect 65102 665618 104546 665854
rect 104782 665618 104866 665854
rect 105102 665618 144546 665854
rect 144782 665618 144866 665854
rect 145102 665618 184546 665854
rect 184782 665618 184866 665854
rect 185102 665618 224546 665854
rect 224782 665618 224866 665854
rect 225102 665618 264546 665854
rect 264782 665618 264866 665854
rect 265102 665618 304546 665854
rect 304782 665618 304866 665854
rect 305102 665618 344546 665854
rect 344782 665618 344866 665854
rect 345102 665618 384546 665854
rect 384782 665618 384866 665854
rect 385102 665618 424546 665854
rect 424782 665618 424866 665854
rect 425102 665618 464546 665854
rect 464782 665618 464866 665854
rect 465102 665618 504546 665854
rect 504782 665618 504866 665854
rect 505102 665618 544546 665854
rect 544782 665618 544866 665854
rect 545102 665618 588222 665854
rect 588458 665618 588542 665854
rect 588778 665618 588810 665854
rect -4886 665586 588810 665618
rect -2966 662454 586890 662486
rect -2966 662218 -2934 662454
rect -2698 662218 -2614 662454
rect -2378 662218 20826 662454
rect 21062 662218 21146 662454
rect 21382 662218 60826 662454
rect 61062 662218 61146 662454
rect 61382 662218 100826 662454
rect 101062 662218 101146 662454
rect 101382 662218 140826 662454
rect 141062 662218 141146 662454
rect 141382 662218 180826 662454
rect 181062 662218 181146 662454
rect 181382 662218 220826 662454
rect 221062 662218 221146 662454
rect 221382 662218 260826 662454
rect 261062 662218 261146 662454
rect 261382 662218 300826 662454
rect 301062 662218 301146 662454
rect 301382 662218 340826 662454
rect 341062 662218 341146 662454
rect 341382 662218 380826 662454
rect 381062 662218 381146 662454
rect 381382 662218 420826 662454
rect 421062 662218 421146 662454
rect 421382 662218 460826 662454
rect 461062 662218 461146 662454
rect 461382 662218 500826 662454
rect 501062 662218 501146 662454
rect 501382 662218 540826 662454
rect 541062 662218 541146 662454
rect 541382 662218 580826 662454
rect 581062 662218 581146 662454
rect 581382 662218 586302 662454
rect 586538 662218 586622 662454
rect 586858 662218 586890 662454
rect -2966 662134 586890 662218
rect -2966 661898 -2934 662134
rect -2698 661898 -2614 662134
rect -2378 661898 20826 662134
rect 21062 661898 21146 662134
rect 21382 661898 60826 662134
rect 61062 661898 61146 662134
rect 61382 661898 100826 662134
rect 101062 661898 101146 662134
rect 101382 661898 140826 662134
rect 141062 661898 141146 662134
rect 141382 661898 180826 662134
rect 181062 661898 181146 662134
rect 181382 661898 220826 662134
rect 221062 661898 221146 662134
rect 221382 661898 260826 662134
rect 261062 661898 261146 662134
rect 261382 661898 300826 662134
rect 301062 661898 301146 662134
rect 301382 661898 340826 662134
rect 341062 661898 341146 662134
rect 341382 661898 380826 662134
rect 381062 661898 381146 662134
rect 381382 661898 420826 662134
rect 421062 661898 421146 662134
rect 421382 661898 460826 662134
rect 461062 661898 461146 662134
rect 461382 661898 500826 662134
rect 501062 661898 501146 662134
rect 501382 661898 540826 662134
rect 541062 661898 541146 662134
rect 541382 661898 580826 662134
rect 581062 661898 581146 662134
rect 581382 661898 586302 662134
rect 586538 661898 586622 662134
rect 586858 661898 586890 662134
rect -2966 661866 586890 661898
rect -8726 653614 592650 653646
rect -8726 653378 -7734 653614
rect -7498 653378 -7414 653614
rect -7178 653378 11986 653614
rect 12222 653378 12306 653614
rect 12542 653378 51986 653614
rect 52222 653378 52306 653614
rect 52542 653378 91986 653614
rect 92222 653378 92306 653614
rect 92542 653378 131986 653614
rect 132222 653378 132306 653614
rect 132542 653378 171986 653614
rect 172222 653378 172306 653614
rect 172542 653378 211986 653614
rect 212222 653378 212306 653614
rect 212542 653378 251986 653614
rect 252222 653378 252306 653614
rect 252542 653378 291986 653614
rect 292222 653378 292306 653614
rect 292542 653378 331986 653614
rect 332222 653378 332306 653614
rect 332542 653378 371986 653614
rect 372222 653378 372306 653614
rect 372542 653378 411986 653614
rect 412222 653378 412306 653614
rect 412542 653378 451986 653614
rect 452222 653378 452306 653614
rect 452542 653378 491986 653614
rect 492222 653378 492306 653614
rect 492542 653378 531986 653614
rect 532222 653378 532306 653614
rect 532542 653378 571986 653614
rect 572222 653378 572306 653614
rect 572542 653378 591102 653614
rect 591338 653378 591422 653614
rect 591658 653378 592650 653614
rect -8726 653294 592650 653378
rect -8726 653058 -7734 653294
rect -7498 653058 -7414 653294
rect -7178 653058 11986 653294
rect 12222 653058 12306 653294
rect 12542 653058 51986 653294
rect 52222 653058 52306 653294
rect 52542 653058 91986 653294
rect 92222 653058 92306 653294
rect 92542 653058 131986 653294
rect 132222 653058 132306 653294
rect 132542 653058 171986 653294
rect 172222 653058 172306 653294
rect 172542 653058 211986 653294
rect 212222 653058 212306 653294
rect 212542 653058 251986 653294
rect 252222 653058 252306 653294
rect 252542 653058 291986 653294
rect 292222 653058 292306 653294
rect 292542 653058 331986 653294
rect 332222 653058 332306 653294
rect 332542 653058 371986 653294
rect 372222 653058 372306 653294
rect 372542 653058 411986 653294
rect 412222 653058 412306 653294
rect 412542 653058 451986 653294
rect 452222 653058 452306 653294
rect 452542 653058 491986 653294
rect 492222 653058 492306 653294
rect 492542 653058 531986 653294
rect 532222 653058 532306 653294
rect 532542 653058 571986 653294
rect 572222 653058 572306 653294
rect 572542 653058 591102 653294
rect 591338 653058 591422 653294
rect 591658 653058 592650 653294
rect -8726 653026 592650 653058
rect -6806 649894 590730 649926
rect -6806 649658 -5814 649894
rect -5578 649658 -5494 649894
rect -5258 649658 8266 649894
rect 8502 649658 8586 649894
rect 8822 649658 48266 649894
rect 48502 649658 48586 649894
rect 48822 649658 88266 649894
rect 88502 649658 88586 649894
rect 88822 649658 128266 649894
rect 128502 649658 128586 649894
rect 128822 649658 168266 649894
rect 168502 649658 168586 649894
rect 168822 649658 208266 649894
rect 208502 649658 208586 649894
rect 208822 649658 248266 649894
rect 248502 649658 248586 649894
rect 248822 649658 288266 649894
rect 288502 649658 288586 649894
rect 288822 649658 328266 649894
rect 328502 649658 328586 649894
rect 328822 649658 368266 649894
rect 368502 649658 368586 649894
rect 368822 649658 408266 649894
rect 408502 649658 408586 649894
rect 408822 649658 448266 649894
rect 448502 649658 448586 649894
rect 448822 649658 488266 649894
rect 488502 649658 488586 649894
rect 488822 649658 528266 649894
rect 528502 649658 528586 649894
rect 528822 649658 568266 649894
rect 568502 649658 568586 649894
rect 568822 649658 589182 649894
rect 589418 649658 589502 649894
rect 589738 649658 590730 649894
rect -6806 649574 590730 649658
rect -6806 649338 -5814 649574
rect -5578 649338 -5494 649574
rect -5258 649338 8266 649574
rect 8502 649338 8586 649574
rect 8822 649338 48266 649574
rect 48502 649338 48586 649574
rect 48822 649338 88266 649574
rect 88502 649338 88586 649574
rect 88822 649338 128266 649574
rect 128502 649338 128586 649574
rect 128822 649338 168266 649574
rect 168502 649338 168586 649574
rect 168822 649338 208266 649574
rect 208502 649338 208586 649574
rect 208822 649338 248266 649574
rect 248502 649338 248586 649574
rect 248822 649338 288266 649574
rect 288502 649338 288586 649574
rect 288822 649338 328266 649574
rect 328502 649338 328586 649574
rect 328822 649338 368266 649574
rect 368502 649338 368586 649574
rect 368822 649338 408266 649574
rect 408502 649338 408586 649574
rect 408822 649338 448266 649574
rect 448502 649338 448586 649574
rect 448822 649338 488266 649574
rect 488502 649338 488586 649574
rect 488822 649338 528266 649574
rect 528502 649338 528586 649574
rect 528822 649338 568266 649574
rect 568502 649338 568586 649574
rect 568822 649338 589182 649574
rect 589418 649338 589502 649574
rect 589738 649338 590730 649574
rect -6806 649306 590730 649338
rect -4886 646174 588810 646206
rect -4886 645938 -3894 646174
rect -3658 645938 -3574 646174
rect -3338 645938 4546 646174
rect 4782 645938 4866 646174
rect 5102 645938 44546 646174
rect 44782 645938 44866 646174
rect 45102 645938 84546 646174
rect 84782 645938 84866 646174
rect 85102 645938 124546 646174
rect 124782 645938 124866 646174
rect 125102 645938 164546 646174
rect 164782 645938 164866 646174
rect 165102 645938 204546 646174
rect 204782 645938 204866 646174
rect 205102 645938 244546 646174
rect 244782 645938 244866 646174
rect 245102 645938 284546 646174
rect 284782 645938 284866 646174
rect 285102 645938 324546 646174
rect 324782 645938 324866 646174
rect 325102 645938 364546 646174
rect 364782 645938 364866 646174
rect 365102 645938 404546 646174
rect 404782 645938 404866 646174
rect 405102 645938 444546 646174
rect 444782 645938 444866 646174
rect 445102 645938 484546 646174
rect 484782 645938 484866 646174
rect 485102 645938 524546 646174
rect 524782 645938 524866 646174
rect 525102 645938 564546 646174
rect 564782 645938 564866 646174
rect 565102 645938 587262 646174
rect 587498 645938 587582 646174
rect 587818 645938 588810 646174
rect -4886 645854 588810 645938
rect -4886 645618 -3894 645854
rect -3658 645618 -3574 645854
rect -3338 645618 4546 645854
rect 4782 645618 4866 645854
rect 5102 645618 44546 645854
rect 44782 645618 44866 645854
rect 45102 645618 84546 645854
rect 84782 645618 84866 645854
rect 85102 645618 124546 645854
rect 124782 645618 124866 645854
rect 125102 645618 164546 645854
rect 164782 645618 164866 645854
rect 165102 645618 204546 645854
rect 204782 645618 204866 645854
rect 205102 645618 244546 645854
rect 244782 645618 244866 645854
rect 245102 645618 284546 645854
rect 284782 645618 284866 645854
rect 285102 645618 324546 645854
rect 324782 645618 324866 645854
rect 325102 645618 364546 645854
rect 364782 645618 364866 645854
rect 365102 645618 404546 645854
rect 404782 645618 404866 645854
rect 405102 645618 444546 645854
rect 444782 645618 444866 645854
rect 445102 645618 484546 645854
rect 484782 645618 484866 645854
rect 485102 645618 524546 645854
rect 524782 645618 524866 645854
rect 525102 645618 564546 645854
rect 564782 645618 564866 645854
rect 565102 645618 587262 645854
rect 587498 645618 587582 645854
rect 587818 645618 588810 645854
rect -4886 645586 588810 645618
rect -2966 642454 586890 642486
rect -2966 642218 -1974 642454
rect -1738 642218 -1654 642454
rect -1418 642218 826 642454
rect 1062 642218 1146 642454
rect 1382 642218 40826 642454
rect 41062 642218 41146 642454
rect 41382 642218 80826 642454
rect 81062 642218 81146 642454
rect 81382 642218 120826 642454
rect 121062 642218 121146 642454
rect 121382 642218 160826 642454
rect 161062 642218 161146 642454
rect 161382 642218 200826 642454
rect 201062 642218 201146 642454
rect 201382 642218 240826 642454
rect 241062 642218 241146 642454
rect 241382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 320826 642454
rect 321062 642218 321146 642454
rect 321382 642218 360826 642454
rect 361062 642218 361146 642454
rect 361382 642218 400826 642454
rect 401062 642218 401146 642454
rect 401382 642218 440826 642454
rect 441062 642218 441146 642454
rect 441382 642218 480826 642454
rect 481062 642218 481146 642454
rect 481382 642218 520826 642454
rect 521062 642218 521146 642454
rect 521382 642218 560826 642454
rect 561062 642218 561146 642454
rect 561382 642218 585342 642454
rect 585578 642218 585662 642454
rect 585898 642218 586890 642454
rect -2966 642134 586890 642218
rect -2966 641898 -1974 642134
rect -1738 641898 -1654 642134
rect -1418 641898 826 642134
rect 1062 641898 1146 642134
rect 1382 641898 40826 642134
rect 41062 641898 41146 642134
rect 41382 641898 80826 642134
rect 81062 641898 81146 642134
rect 81382 641898 120826 642134
rect 121062 641898 121146 642134
rect 121382 641898 160826 642134
rect 161062 641898 161146 642134
rect 161382 641898 200826 642134
rect 201062 641898 201146 642134
rect 201382 641898 240826 642134
rect 241062 641898 241146 642134
rect 241382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 320826 642134
rect 321062 641898 321146 642134
rect 321382 641898 360826 642134
rect 361062 641898 361146 642134
rect 361382 641898 400826 642134
rect 401062 641898 401146 642134
rect 401382 641898 440826 642134
rect 441062 641898 441146 642134
rect 441382 641898 480826 642134
rect 481062 641898 481146 642134
rect 481382 641898 520826 642134
rect 521062 641898 521146 642134
rect 521382 641898 560826 642134
rect 561062 641898 561146 642134
rect 561382 641898 585342 642134
rect 585578 641898 585662 642134
rect 585898 641898 586890 642134
rect -2966 641866 586890 641898
rect -8726 633614 592650 633646
rect -8726 633378 -8694 633614
rect -8458 633378 -8374 633614
rect -8138 633378 31986 633614
rect 32222 633378 32306 633614
rect 32542 633378 71986 633614
rect 72222 633378 72306 633614
rect 72542 633378 111986 633614
rect 112222 633378 112306 633614
rect 112542 633378 151986 633614
rect 152222 633378 152306 633614
rect 152542 633378 191986 633614
rect 192222 633378 192306 633614
rect 192542 633378 231986 633614
rect 232222 633378 232306 633614
rect 232542 633378 271986 633614
rect 272222 633378 272306 633614
rect 272542 633378 311986 633614
rect 312222 633378 312306 633614
rect 312542 633378 351986 633614
rect 352222 633378 352306 633614
rect 352542 633378 391986 633614
rect 392222 633378 392306 633614
rect 392542 633378 431986 633614
rect 432222 633378 432306 633614
rect 432542 633378 471986 633614
rect 472222 633378 472306 633614
rect 472542 633378 511986 633614
rect 512222 633378 512306 633614
rect 512542 633378 551986 633614
rect 552222 633378 552306 633614
rect 552542 633378 592062 633614
rect 592298 633378 592382 633614
rect 592618 633378 592650 633614
rect -8726 633294 592650 633378
rect -8726 633058 -8694 633294
rect -8458 633058 -8374 633294
rect -8138 633058 31986 633294
rect 32222 633058 32306 633294
rect 32542 633058 71986 633294
rect 72222 633058 72306 633294
rect 72542 633058 111986 633294
rect 112222 633058 112306 633294
rect 112542 633058 151986 633294
rect 152222 633058 152306 633294
rect 152542 633058 191986 633294
rect 192222 633058 192306 633294
rect 192542 633058 231986 633294
rect 232222 633058 232306 633294
rect 232542 633058 271986 633294
rect 272222 633058 272306 633294
rect 272542 633058 311986 633294
rect 312222 633058 312306 633294
rect 312542 633058 351986 633294
rect 352222 633058 352306 633294
rect 352542 633058 391986 633294
rect 392222 633058 392306 633294
rect 392542 633058 431986 633294
rect 432222 633058 432306 633294
rect 432542 633058 471986 633294
rect 472222 633058 472306 633294
rect 472542 633058 511986 633294
rect 512222 633058 512306 633294
rect 512542 633058 551986 633294
rect 552222 633058 552306 633294
rect 552542 633058 592062 633294
rect 592298 633058 592382 633294
rect 592618 633058 592650 633294
rect -8726 633026 592650 633058
rect -6806 629894 590730 629926
rect -6806 629658 -6774 629894
rect -6538 629658 -6454 629894
rect -6218 629658 28266 629894
rect 28502 629658 28586 629894
rect 28822 629658 68266 629894
rect 68502 629658 68586 629894
rect 68822 629658 108266 629894
rect 108502 629658 108586 629894
rect 108822 629658 148266 629894
rect 148502 629658 148586 629894
rect 148822 629658 188266 629894
rect 188502 629658 188586 629894
rect 188822 629658 228266 629894
rect 228502 629658 228586 629894
rect 228822 629658 268266 629894
rect 268502 629658 268586 629894
rect 268822 629658 308266 629894
rect 308502 629658 308586 629894
rect 308822 629658 348266 629894
rect 348502 629658 348586 629894
rect 348822 629658 388266 629894
rect 388502 629658 388586 629894
rect 388822 629658 428266 629894
rect 428502 629658 428586 629894
rect 428822 629658 468266 629894
rect 468502 629658 468586 629894
rect 468822 629658 508266 629894
rect 508502 629658 508586 629894
rect 508822 629658 548266 629894
rect 548502 629658 548586 629894
rect 548822 629658 590142 629894
rect 590378 629658 590462 629894
rect 590698 629658 590730 629894
rect -6806 629574 590730 629658
rect -6806 629338 -6774 629574
rect -6538 629338 -6454 629574
rect -6218 629338 28266 629574
rect 28502 629338 28586 629574
rect 28822 629338 68266 629574
rect 68502 629338 68586 629574
rect 68822 629338 108266 629574
rect 108502 629338 108586 629574
rect 108822 629338 148266 629574
rect 148502 629338 148586 629574
rect 148822 629338 188266 629574
rect 188502 629338 188586 629574
rect 188822 629338 228266 629574
rect 228502 629338 228586 629574
rect 228822 629338 268266 629574
rect 268502 629338 268586 629574
rect 268822 629338 308266 629574
rect 308502 629338 308586 629574
rect 308822 629338 348266 629574
rect 348502 629338 348586 629574
rect 348822 629338 388266 629574
rect 388502 629338 388586 629574
rect 388822 629338 428266 629574
rect 428502 629338 428586 629574
rect 428822 629338 468266 629574
rect 468502 629338 468586 629574
rect 468822 629338 508266 629574
rect 508502 629338 508586 629574
rect 508822 629338 548266 629574
rect 548502 629338 548586 629574
rect 548822 629338 590142 629574
rect 590378 629338 590462 629574
rect 590698 629338 590730 629574
rect -6806 629306 590730 629338
rect -4886 626174 588810 626206
rect -4886 625938 -4854 626174
rect -4618 625938 -4534 626174
rect -4298 625938 24546 626174
rect 24782 625938 24866 626174
rect 25102 625938 64546 626174
rect 64782 625938 64866 626174
rect 65102 625938 104546 626174
rect 104782 625938 104866 626174
rect 105102 625938 144546 626174
rect 144782 625938 144866 626174
rect 145102 625938 184546 626174
rect 184782 625938 184866 626174
rect 185102 625938 224546 626174
rect 224782 625938 224866 626174
rect 225102 625938 264546 626174
rect 264782 625938 264866 626174
rect 265102 625938 304546 626174
rect 304782 625938 304866 626174
rect 305102 625938 344546 626174
rect 344782 625938 344866 626174
rect 345102 625938 384546 626174
rect 384782 625938 384866 626174
rect 385102 625938 424546 626174
rect 424782 625938 424866 626174
rect 425102 625938 464546 626174
rect 464782 625938 464866 626174
rect 465102 625938 504546 626174
rect 504782 625938 504866 626174
rect 505102 625938 544546 626174
rect 544782 625938 544866 626174
rect 545102 625938 588222 626174
rect 588458 625938 588542 626174
rect 588778 625938 588810 626174
rect -4886 625854 588810 625938
rect -4886 625618 -4854 625854
rect -4618 625618 -4534 625854
rect -4298 625618 24546 625854
rect 24782 625618 24866 625854
rect 25102 625618 64546 625854
rect 64782 625618 64866 625854
rect 65102 625618 104546 625854
rect 104782 625618 104866 625854
rect 105102 625618 144546 625854
rect 144782 625618 144866 625854
rect 145102 625618 184546 625854
rect 184782 625618 184866 625854
rect 185102 625618 224546 625854
rect 224782 625618 224866 625854
rect 225102 625618 264546 625854
rect 264782 625618 264866 625854
rect 265102 625618 304546 625854
rect 304782 625618 304866 625854
rect 305102 625618 344546 625854
rect 344782 625618 344866 625854
rect 345102 625618 384546 625854
rect 384782 625618 384866 625854
rect 385102 625618 424546 625854
rect 424782 625618 424866 625854
rect 425102 625618 464546 625854
rect 464782 625618 464866 625854
rect 465102 625618 504546 625854
rect 504782 625618 504866 625854
rect 505102 625618 544546 625854
rect 544782 625618 544866 625854
rect 545102 625618 588222 625854
rect 588458 625618 588542 625854
rect 588778 625618 588810 625854
rect -4886 625586 588810 625618
rect -2966 622454 586890 622486
rect -2966 622218 -2934 622454
rect -2698 622218 -2614 622454
rect -2378 622218 20826 622454
rect 21062 622218 21146 622454
rect 21382 622218 60826 622454
rect 61062 622218 61146 622454
rect 61382 622218 100826 622454
rect 101062 622218 101146 622454
rect 101382 622218 140826 622454
rect 141062 622218 141146 622454
rect 141382 622218 180826 622454
rect 181062 622218 181146 622454
rect 181382 622218 220826 622454
rect 221062 622218 221146 622454
rect 221382 622218 260826 622454
rect 261062 622218 261146 622454
rect 261382 622218 300826 622454
rect 301062 622218 301146 622454
rect 301382 622218 340826 622454
rect 341062 622218 341146 622454
rect 341382 622218 380826 622454
rect 381062 622218 381146 622454
rect 381382 622218 420826 622454
rect 421062 622218 421146 622454
rect 421382 622218 460826 622454
rect 461062 622218 461146 622454
rect 461382 622218 500826 622454
rect 501062 622218 501146 622454
rect 501382 622218 540826 622454
rect 541062 622218 541146 622454
rect 541382 622218 580826 622454
rect 581062 622218 581146 622454
rect 581382 622218 586302 622454
rect 586538 622218 586622 622454
rect 586858 622218 586890 622454
rect -2966 622134 586890 622218
rect -2966 621898 -2934 622134
rect -2698 621898 -2614 622134
rect -2378 621898 20826 622134
rect 21062 621898 21146 622134
rect 21382 621898 60826 622134
rect 61062 621898 61146 622134
rect 61382 621898 100826 622134
rect 101062 621898 101146 622134
rect 101382 621898 140826 622134
rect 141062 621898 141146 622134
rect 141382 621898 180826 622134
rect 181062 621898 181146 622134
rect 181382 621898 220826 622134
rect 221062 621898 221146 622134
rect 221382 621898 260826 622134
rect 261062 621898 261146 622134
rect 261382 621898 300826 622134
rect 301062 621898 301146 622134
rect 301382 621898 340826 622134
rect 341062 621898 341146 622134
rect 341382 621898 380826 622134
rect 381062 621898 381146 622134
rect 381382 621898 420826 622134
rect 421062 621898 421146 622134
rect 421382 621898 460826 622134
rect 461062 621898 461146 622134
rect 461382 621898 500826 622134
rect 501062 621898 501146 622134
rect 501382 621898 540826 622134
rect 541062 621898 541146 622134
rect 541382 621898 580826 622134
rect 581062 621898 581146 622134
rect 581382 621898 586302 622134
rect 586538 621898 586622 622134
rect 586858 621898 586890 622134
rect -2966 621866 586890 621898
rect -8726 613614 592650 613646
rect -8726 613378 -7734 613614
rect -7498 613378 -7414 613614
rect -7178 613378 11986 613614
rect 12222 613378 12306 613614
rect 12542 613378 51986 613614
rect 52222 613378 52306 613614
rect 52542 613378 91986 613614
rect 92222 613378 92306 613614
rect 92542 613378 131986 613614
rect 132222 613378 132306 613614
rect 132542 613378 171986 613614
rect 172222 613378 172306 613614
rect 172542 613378 211986 613614
rect 212222 613378 212306 613614
rect 212542 613378 251986 613614
rect 252222 613378 252306 613614
rect 252542 613378 291986 613614
rect 292222 613378 292306 613614
rect 292542 613378 331986 613614
rect 332222 613378 332306 613614
rect 332542 613378 371986 613614
rect 372222 613378 372306 613614
rect 372542 613378 411986 613614
rect 412222 613378 412306 613614
rect 412542 613378 451986 613614
rect 452222 613378 452306 613614
rect 452542 613378 491986 613614
rect 492222 613378 492306 613614
rect 492542 613378 531986 613614
rect 532222 613378 532306 613614
rect 532542 613378 571986 613614
rect 572222 613378 572306 613614
rect 572542 613378 591102 613614
rect 591338 613378 591422 613614
rect 591658 613378 592650 613614
rect -8726 613294 592650 613378
rect -8726 613058 -7734 613294
rect -7498 613058 -7414 613294
rect -7178 613058 11986 613294
rect 12222 613058 12306 613294
rect 12542 613058 51986 613294
rect 52222 613058 52306 613294
rect 52542 613058 91986 613294
rect 92222 613058 92306 613294
rect 92542 613058 131986 613294
rect 132222 613058 132306 613294
rect 132542 613058 171986 613294
rect 172222 613058 172306 613294
rect 172542 613058 211986 613294
rect 212222 613058 212306 613294
rect 212542 613058 251986 613294
rect 252222 613058 252306 613294
rect 252542 613058 291986 613294
rect 292222 613058 292306 613294
rect 292542 613058 331986 613294
rect 332222 613058 332306 613294
rect 332542 613058 371986 613294
rect 372222 613058 372306 613294
rect 372542 613058 411986 613294
rect 412222 613058 412306 613294
rect 412542 613058 451986 613294
rect 452222 613058 452306 613294
rect 452542 613058 491986 613294
rect 492222 613058 492306 613294
rect 492542 613058 531986 613294
rect 532222 613058 532306 613294
rect 532542 613058 571986 613294
rect 572222 613058 572306 613294
rect 572542 613058 591102 613294
rect 591338 613058 591422 613294
rect 591658 613058 592650 613294
rect -8726 613026 592650 613058
rect -6806 609894 590730 609926
rect -6806 609658 -5814 609894
rect -5578 609658 -5494 609894
rect -5258 609658 8266 609894
rect 8502 609658 8586 609894
rect 8822 609658 48266 609894
rect 48502 609658 48586 609894
rect 48822 609658 88266 609894
rect 88502 609658 88586 609894
rect 88822 609658 128266 609894
rect 128502 609658 128586 609894
rect 128822 609658 168266 609894
rect 168502 609658 168586 609894
rect 168822 609658 208266 609894
rect 208502 609658 208586 609894
rect 208822 609658 248266 609894
rect 248502 609658 248586 609894
rect 248822 609658 288266 609894
rect 288502 609658 288586 609894
rect 288822 609658 328266 609894
rect 328502 609658 328586 609894
rect 328822 609658 368266 609894
rect 368502 609658 368586 609894
rect 368822 609658 408266 609894
rect 408502 609658 408586 609894
rect 408822 609658 448266 609894
rect 448502 609658 448586 609894
rect 448822 609658 488266 609894
rect 488502 609658 488586 609894
rect 488822 609658 528266 609894
rect 528502 609658 528586 609894
rect 528822 609658 568266 609894
rect 568502 609658 568586 609894
rect 568822 609658 589182 609894
rect 589418 609658 589502 609894
rect 589738 609658 590730 609894
rect -6806 609574 590730 609658
rect -6806 609338 -5814 609574
rect -5578 609338 -5494 609574
rect -5258 609338 8266 609574
rect 8502 609338 8586 609574
rect 8822 609338 48266 609574
rect 48502 609338 48586 609574
rect 48822 609338 88266 609574
rect 88502 609338 88586 609574
rect 88822 609338 128266 609574
rect 128502 609338 128586 609574
rect 128822 609338 168266 609574
rect 168502 609338 168586 609574
rect 168822 609338 208266 609574
rect 208502 609338 208586 609574
rect 208822 609338 248266 609574
rect 248502 609338 248586 609574
rect 248822 609338 288266 609574
rect 288502 609338 288586 609574
rect 288822 609338 328266 609574
rect 328502 609338 328586 609574
rect 328822 609338 368266 609574
rect 368502 609338 368586 609574
rect 368822 609338 408266 609574
rect 408502 609338 408586 609574
rect 408822 609338 448266 609574
rect 448502 609338 448586 609574
rect 448822 609338 488266 609574
rect 488502 609338 488586 609574
rect 488822 609338 528266 609574
rect 528502 609338 528586 609574
rect 528822 609338 568266 609574
rect 568502 609338 568586 609574
rect 568822 609338 589182 609574
rect 589418 609338 589502 609574
rect 589738 609338 590730 609574
rect -6806 609306 590730 609338
rect -4886 606174 588810 606206
rect -4886 605938 -3894 606174
rect -3658 605938 -3574 606174
rect -3338 605938 4546 606174
rect 4782 605938 4866 606174
rect 5102 605938 44546 606174
rect 44782 605938 44866 606174
rect 45102 605938 84546 606174
rect 84782 605938 84866 606174
rect 85102 605938 124546 606174
rect 124782 605938 124866 606174
rect 125102 605938 164546 606174
rect 164782 605938 164866 606174
rect 165102 605938 204546 606174
rect 204782 605938 204866 606174
rect 205102 605938 244546 606174
rect 244782 605938 244866 606174
rect 245102 605938 284546 606174
rect 284782 605938 284866 606174
rect 285102 605938 324546 606174
rect 324782 605938 324866 606174
rect 325102 605938 364546 606174
rect 364782 605938 364866 606174
rect 365102 605938 404546 606174
rect 404782 605938 404866 606174
rect 405102 605938 444546 606174
rect 444782 605938 444866 606174
rect 445102 605938 484546 606174
rect 484782 605938 484866 606174
rect 485102 605938 524546 606174
rect 524782 605938 524866 606174
rect 525102 605938 564546 606174
rect 564782 605938 564866 606174
rect 565102 605938 587262 606174
rect 587498 605938 587582 606174
rect 587818 605938 588810 606174
rect -4886 605854 588810 605938
rect -4886 605618 -3894 605854
rect -3658 605618 -3574 605854
rect -3338 605618 4546 605854
rect 4782 605618 4866 605854
rect 5102 605618 44546 605854
rect 44782 605618 44866 605854
rect 45102 605618 84546 605854
rect 84782 605618 84866 605854
rect 85102 605618 124546 605854
rect 124782 605618 124866 605854
rect 125102 605618 164546 605854
rect 164782 605618 164866 605854
rect 165102 605618 204546 605854
rect 204782 605618 204866 605854
rect 205102 605618 244546 605854
rect 244782 605618 244866 605854
rect 245102 605618 284546 605854
rect 284782 605618 284866 605854
rect 285102 605618 324546 605854
rect 324782 605618 324866 605854
rect 325102 605618 364546 605854
rect 364782 605618 364866 605854
rect 365102 605618 404546 605854
rect 404782 605618 404866 605854
rect 405102 605618 444546 605854
rect 444782 605618 444866 605854
rect 445102 605618 484546 605854
rect 484782 605618 484866 605854
rect 485102 605618 524546 605854
rect 524782 605618 524866 605854
rect 525102 605618 564546 605854
rect 564782 605618 564866 605854
rect 565102 605618 587262 605854
rect 587498 605618 587582 605854
rect 587818 605618 588810 605854
rect -4886 605586 588810 605618
rect -2966 602454 586890 602486
rect -2966 602218 -1974 602454
rect -1738 602218 -1654 602454
rect -1418 602218 826 602454
rect 1062 602218 1146 602454
rect 1382 602218 40826 602454
rect 41062 602218 41146 602454
rect 41382 602218 80826 602454
rect 81062 602218 81146 602454
rect 81382 602218 120826 602454
rect 121062 602218 121146 602454
rect 121382 602218 160826 602454
rect 161062 602218 161146 602454
rect 161382 602218 200826 602454
rect 201062 602218 201146 602454
rect 201382 602218 240826 602454
rect 241062 602218 241146 602454
rect 241382 602218 280826 602454
rect 281062 602218 281146 602454
rect 281382 602218 320826 602454
rect 321062 602218 321146 602454
rect 321382 602218 360826 602454
rect 361062 602218 361146 602454
rect 361382 602218 400826 602454
rect 401062 602218 401146 602454
rect 401382 602218 440826 602454
rect 441062 602218 441146 602454
rect 441382 602218 480826 602454
rect 481062 602218 481146 602454
rect 481382 602218 520826 602454
rect 521062 602218 521146 602454
rect 521382 602218 560826 602454
rect 561062 602218 561146 602454
rect 561382 602218 585342 602454
rect 585578 602218 585662 602454
rect 585898 602218 586890 602454
rect -2966 602134 586890 602218
rect -2966 601898 -1974 602134
rect -1738 601898 -1654 602134
rect -1418 601898 826 602134
rect 1062 601898 1146 602134
rect 1382 601898 40826 602134
rect 41062 601898 41146 602134
rect 41382 601898 80826 602134
rect 81062 601898 81146 602134
rect 81382 601898 120826 602134
rect 121062 601898 121146 602134
rect 121382 601898 160826 602134
rect 161062 601898 161146 602134
rect 161382 601898 200826 602134
rect 201062 601898 201146 602134
rect 201382 601898 240826 602134
rect 241062 601898 241146 602134
rect 241382 601898 280826 602134
rect 281062 601898 281146 602134
rect 281382 601898 320826 602134
rect 321062 601898 321146 602134
rect 321382 601898 360826 602134
rect 361062 601898 361146 602134
rect 361382 601898 400826 602134
rect 401062 601898 401146 602134
rect 401382 601898 440826 602134
rect 441062 601898 441146 602134
rect 441382 601898 480826 602134
rect 481062 601898 481146 602134
rect 481382 601898 520826 602134
rect 521062 601898 521146 602134
rect 521382 601898 560826 602134
rect 561062 601898 561146 602134
rect 561382 601898 585342 602134
rect 585578 601898 585662 602134
rect 585898 601898 586890 602134
rect -2966 601866 586890 601898
rect -8726 593614 592650 593646
rect -8726 593378 -8694 593614
rect -8458 593378 -8374 593614
rect -8138 593378 31986 593614
rect 32222 593378 32306 593614
rect 32542 593378 71986 593614
rect 72222 593378 72306 593614
rect 72542 593378 111986 593614
rect 112222 593378 112306 593614
rect 112542 593378 151986 593614
rect 152222 593378 152306 593614
rect 152542 593378 191986 593614
rect 192222 593378 192306 593614
rect 192542 593378 231986 593614
rect 232222 593378 232306 593614
rect 232542 593378 271986 593614
rect 272222 593378 272306 593614
rect 272542 593378 311986 593614
rect 312222 593378 312306 593614
rect 312542 593378 351986 593614
rect 352222 593378 352306 593614
rect 352542 593378 391986 593614
rect 392222 593378 392306 593614
rect 392542 593378 431986 593614
rect 432222 593378 432306 593614
rect 432542 593378 471986 593614
rect 472222 593378 472306 593614
rect 472542 593378 511986 593614
rect 512222 593378 512306 593614
rect 512542 593378 551986 593614
rect 552222 593378 552306 593614
rect 552542 593378 592062 593614
rect 592298 593378 592382 593614
rect 592618 593378 592650 593614
rect -8726 593294 592650 593378
rect -8726 593058 -8694 593294
rect -8458 593058 -8374 593294
rect -8138 593058 31986 593294
rect 32222 593058 32306 593294
rect 32542 593058 71986 593294
rect 72222 593058 72306 593294
rect 72542 593058 111986 593294
rect 112222 593058 112306 593294
rect 112542 593058 151986 593294
rect 152222 593058 152306 593294
rect 152542 593058 191986 593294
rect 192222 593058 192306 593294
rect 192542 593058 231986 593294
rect 232222 593058 232306 593294
rect 232542 593058 271986 593294
rect 272222 593058 272306 593294
rect 272542 593058 311986 593294
rect 312222 593058 312306 593294
rect 312542 593058 351986 593294
rect 352222 593058 352306 593294
rect 352542 593058 391986 593294
rect 392222 593058 392306 593294
rect 392542 593058 431986 593294
rect 432222 593058 432306 593294
rect 432542 593058 471986 593294
rect 472222 593058 472306 593294
rect 472542 593058 511986 593294
rect 512222 593058 512306 593294
rect 512542 593058 551986 593294
rect 552222 593058 552306 593294
rect 552542 593058 592062 593294
rect 592298 593058 592382 593294
rect 592618 593058 592650 593294
rect -8726 593026 592650 593058
rect -6806 589894 590730 589926
rect -6806 589658 -6774 589894
rect -6538 589658 -6454 589894
rect -6218 589658 28266 589894
rect 28502 589658 28586 589894
rect 28822 589658 68266 589894
rect 68502 589658 68586 589894
rect 68822 589658 108266 589894
rect 108502 589658 108586 589894
rect 108822 589658 148266 589894
rect 148502 589658 148586 589894
rect 148822 589658 188266 589894
rect 188502 589658 188586 589894
rect 188822 589658 228266 589894
rect 228502 589658 228586 589894
rect 228822 589658 268266 589894
rect 268502 589658 268586 589894
rect 268822 589658 308266 589894
rect 308502 589658 308586 589894
rect 308822 589658 348266 589894
rect 348502 589658 348586 589894
rect 348822 589658 388266 589894
rect 388502 589658 388586 589894
rect 388822 589658 428266 589894
rect 428502 589658 428586 589894
rect 428822 589658 468266 589894
rect 468502 589658 468586 589894
rect 468822 589658 508266 589894
rect 508502 589658 508586 589894
rect 508822 589658 548266 589894
rect 548502 589658 548586 589894
rect 548822 589658 590142 589894
rect 590378 589658 590462 589894
rect 590698 589658 590730 589894
rect -6806 589574 590730 589658
rect -6806 589338 -6774 589574
rect -6538 589338 -6454 589574
rect -6218 589338 28266 589574
rect 28502 589338 28586 589574
rect 28822 589338 68266 589574
rect 68502 589338 68586 589574
rect 68822 589338 108266 589574
rect 108502 589338 108586 589574
rect 108822 589338 148266 589574
rect 148502 589338 148586 589574
rect 148822 589338 188266 589574
rect 188502 589338 188586 589574
rect 188822 589338 228266 589574
rect 228502 589338 228586 589574
rect 228822 589338 268266 589574
rect 268502 589338 268586 589574
rect 268822 589338 308266 589574
rect 308502 589338 308586 589574
rect 308822 589338 348266 589574
rect 348502 589338 348586 589574
rect 348822 589338 388266 589574
rect 388502 589338 388586 589574
rect 388822 589338 428266 589574
rect 428502 589338 428586 589574
rect 428822 589338 468266 589574
rect 468502 589338 468586 589574
rect 468822 589338 508266 589574
rect 508502 589338 508586 589574
rect 508822 589338 548266 589574
rect 548502 589338 548586 589574
rect 548822 589338 590142 589574
rect 590378 589338 590462 589574
rect 590698 589338 590730 589574
rect -6806 589306 590730 589338
rect -4886 586174 588810 586206
rect -4886 585938 -4854 586174
rect -4618 585938 -4534 586174
rect -4298 585938 24546 586174
rect 24782 585938 24866 586174
rect 25102 585938 64546 586174
rect 64782 585938 64866 586174
rect 65102 585938 104546 586174
rect 104782 585938 104866 586174
rect 105102 585938 144546 586174
rect 144782 585938 144866 586174
rect 145102 585938 184546 586174
rect 184782 585938 184866 586174
rect 185102 585938 224546 586174
rect 224782 585938 224866 586174
rect 225102 585938 264546 586174
rect 264782 585938 264866 586174
rect 265102 585938 304546 586174
rect 304782 585938 304866 586174
rect 305102 585938 344546 586174
rect 344782 585938 344866 586174
rect 345102 585938 384546 586174
rect 384782 585938 384866 586174
rect 385102 585938 424546 586174
rect 424782 585938 424866 586174
rect 425102 585938 464546 586174
rect 464782 585938 464866 586174
rect 465102 585938 504546 586174
rect 504782 585938 504866 586174
rect 505102 585938 544546 586174
rect 544782 585938 544866 586174
rect 545102 585938 588222 586174
rect 588458 585938 588542 586174
rect 588778 585938 588810 586174
rect -4886 585854 588810 585938
rect -4886 585618 -4854 585854
rect -4618 585618 -4534 585854
rect -4298 585618 24546 585854
rect 24782 585618 24866 585854
rect 25102 585618 64546 585854
rect 64782 585618 64866 585854
rect 65102 585618 104546 585854
rect 104782 585618 104866 585854
rect 105102 585618 144546 585854
rect 144782 585618 144866 585854
rect 145102 585618 184546 585854
rect 184782 585618 184866 585854
rect 185102 585618 224546 585854
rect 224782 585618 224866 585854
rect 225102 585618 264546 585854
rect 264782 585618 264866 585854
rect 265102 585618 304546 585854
rect 304782 585618 304866 585854
rect 305102 585618 344546 585854
rect 344782 585618 344866 585854
rect 345102 585618 384546 585854
rect 384782 585618 384866 585854
rect 385102 585618 424546 585854
rect 424782 585618 424866 585854
rect 425102 585618 464546 585854
rect 464782 585618 464866 585854
rect 465102 585618 504546 585854
rect 504782 585618 504866 585854
rect 505102 585618 544546 585854
rect 544782 585618 544866 585854
rect 545102 585618 588222 585854
rect 588458 585618 588542 585854
rect 588778 585618 588810 585854
rect -4886 585586 588810 585618
rect -2966 582454 586890 582486
rect -2966 582218 -2934 582454
rect -2698 582218 -2614 582454
rect -2378 582218 20826 582454
rect 21062 582218 21146 582454
rect 21382 582218 60826 582454
rect 61062 582218 61146 582454
rect 61382 582218 100826 582454
rect 101062 582218 101146 582454
rect 101382 582218 140826 582454
rect 141062 582218 141146 582454
rect 141382 582218 180826 582454
rect 181062 582218 181146 582454
rect 181382 582218 220826 582454
rect 221062 582218 221146 582454
rect 221382 582218 260826 582454
rect 261062 582218 261146 582454
rect 261382 582218 300826 582454
rect 301062 582218 301146 582454
rect 301382 582218 340826 582454
rect 341062 582218 341146 582454
rect 341382 582218 380826 582454
rect 381062 582218 381146 582454
rect 381382 582218 420826 582454
rect 421062 582218 421146 582454
rect 421382 582218 460826 582454
rect 461062 582218 461146 582454
rect 461382 582218 500826 582454
rect 501062 582218 501146 582454
rect 501382 582218 540826 582454
rect 541062 582218 541146 582454
rect 541382 582218 580826 582454
rect 581062 582218 581146 582454
rect 581382 582218 586302 582454
rect 586538 582218 586622 582454
rect 586858 582218 586890 582454
rect -2966 582134 586890 582218
rect -2966 581898 -2934 582134
rect -2698 581898 -2614 582134
rect -2378 581898 20826 582134
rect 21062 581898 21146 582134
rect 21382 581898 60826 582134
rect 61062 581898 61146 582134
rect 61382 581898 100826 582134
rect 101062 581898 101146 582134
rect 101382 581898 140826 582134
rect 141062 581898 141146 582134
rect 141382 581898 180826 582134
rect 181062 581898 181146 582134
rect 181382 581898 220826 582134
rect 221062 581898 221146 582134
rect 221382 581898 260826 582134
rect 261062 581898 261146 582134
rect 261382 581898 300826 582134
rect 301062 581898 301146 582134
rect 301382 581898 340826 582134
rect 341062 581898 341146 582134
rect 341382 581898 380826 582134
rect 381062 581898 381146 582134
rect 381382 581898 420826 582134
rect 421062 581898 421146 582134
rect 421382 581898 460826 582134
rect 461062 581898 461146 582134
rect 461382 581898 500826 582134
rect 501062 581898 501146 582134
rect 501382 581898 540826 582134
rect 541062 581898 541146 582134
rect 541382 581898 580826 582134
rect 581062 581898 581146 582134
rect 581382 581898 586302 582134
rect 586538 581898 586622 582134
rect 586858 581898 586890 582134
rect -2966 581866 586890 581898
rect -8726 573614 592650 573646
rect -8726 573378 -7734 573614
rect -7498 573378 -7414 573614
rect -7178 573378 11986 573614
rect 12222 573378 12306 573614
rect 12542 573378 51986 573614
rect 52222 573378 52306 573614
rect 52542 573378 91986 573614
rect 92222 573378 92306 573614
rect 92542 573378 131986 573614
rect 132222 573378 132306 573614
rect 132542 573378 171986 573614
rect 172222 573378 172306 573614
rect 172542 573378 211986 573614
rect 212222 573378 212306 573614
rect 212542 573378 251986 573614
rect 252222 573378 252306 573614
rect 252542 573378 291986 573614
rect 292222 573378 292306 573614
rect 292542 573378 331986 573614
rect 332222 573378 332306 573614
rect 332542 573378 371986 573614
rect 372222 573378 372306 573614
rect 372542 573378 411986 573614
rect 412222 573378 412306 573614
rect 412542 573378 451986 573614
rect 452222 573378 452306 573614
rect 452542 573378 491986 573614
rect 492222 573378 492306 573614
rect 492542 573378 531986 573614
rect 532222 573378 532306 573614
rect 532542 573378 571986 573614
rect 572222 573378 572306 573614
rect 572542 573378 591102 573614
rect 591338 573378 591422 573614
rect 591658 573378 592650 573614
rect -8726 573294 592650 573378
rect -8726 573058 -7734 573294
rect -7498 573058 -7414 573294
rect -7178 573058 11986 573294
rect 12222 573058 12306 573294
rect 12542 573058 51986 573294
rect 52222 573058 52306 573294
rect 52542 573058 91986 573294
rect 92222 573058 92306 573294
rect 92542 573058 131986 573294
rect 132222 573058 132306 573294
rect 132542 573058 171986 573294
rect 172222 573058 172306 573294
rect 172542 573058 211986 573294
rect 212222 573058 212306 573294
rect 212542 573058 251986 573294
rect 252222 573058 252306 573294
rect 252542 573058 291986 573294
rect 292222 573058 292306 573294
rect 292542 573058 331986 573294
rect 332222 573058 332306 573294
rect 332542 573058 371986 573294
rect 372222 573058 372306 573294
rect 372542 573058 411986 573294
rect 412222 573058 412306 573294
rect 412542 573058 451986 573294
rect 452222 573058 452306 573294
rect 452542 573058 491986 573294
rect 492222 573058 492306 573294
rect 492542 573058 531986 573294
rect 532222 573058 532306 573294
rect 532542 573058 571986 573294
rect 572222 573058 572306 573294
rect 572542 573058 591102 573294
rect 591338 573058 591422 573294
rect 591658 573058 592650 573294
rect -8726 573026 592650 573058
rect -6806 569894 590730 569926
rect -6806 569658 -5814 569894
rect -5578 569658 -5494 569894
rect -5258 569658 8266 569894
rect 8502 569658 8586 569894
rect 8822 569658 48266 569894
rect 48502 569658 48586 569894
rect 48822 569658 88266 569894
rect 88502 569658 88586 569894
rect 88822 569658 128266 569894
rect 128502 569658 128586 569894
rect 128822 569658 168266 569894
rect 168502 569658 168586 569894
rect 168822 569658 208266 569894
rect 208502 569658 208586 569894
rect 208822 569658 248266 569894
rect 248502 569658 248586 569894
rect 248822 569658 288266 569894
rect 288502 569658 288586 569894
rect 288822 569658 328266 569894
rect 328502 569658 328586 569894
rect 328822 569658 368266 569894
rect 368502 569658 368586 569894
rect 368822 569658 408266 569894
rect 408502 569658 408586 569894
rect 408822 569658 448266 569894
rect 448502 569658 448586 569894
rect 448822 569658 488266 569894
rect 488502 569658 488586 569894
rect 488822 569658 528266 569894
rect 528502 569658 528586 569894
rect 528822 569658 568266 569894
rect 568502 569658 568586 569894
rect 568822 569658 589182 569894
rect 589418 569658 589502 569894
rect 589738 569658 590730 569894
rect -6806 569574 590730 569658
rect -6806 569338 -5814 569574
rect -5578 569338 -5494 569574
rect -5258 569338 8266 569574
rect 8502 569338 8586 569574
rect 8822 569338 48266 569574
rect 48502 569338 48586 569574
rect 48822 569338 88266 569574
rect 88502 569338 88586 569574
rect 88822 569338 128266 569574
rect 128502 569338 128586 569574
rect 128822 569338 168266 569574
rect 168502 569338 168586 569574
rect 168822 569338 208266 569574
rect 208502 569338 208586 569574
rect 208822 569338 248266 569574
rect 248502 569338 248586 569574
rect 248822 569338 288266 569574
rect 288502 569338 288586 569574
rect 288822 569338 328266 569574
rect 328502 569338 328586 569574
rect 328822 569338 368266 569574
rect 368502 569338 368586 569574
rect 368822 569338 408266 569574
rect 408502 569338 408586 569574
rect 408822 569338 448266 569574
rect 448502 569338 448586 569574
rect 448822 569338 488266 569574
rect 488502 569338 488586 569574
rect 488822 569338 528266 569574
rect 528502 569338 528586 569574
rect 528822 569338 568266 569574
rect 568502 569338 568586 569574
rect 568822 569338 589182 569574
rect 589418 569338 589502 569574
rect 589738 569338 590730 569574
rect -6806 569306 590730 569338
rect -4886 566174 588810 566206
rect -4886 565938 -3894 566174
rect -3658 565938 -3574 566174
rect -3338 565938 4546 566174
rect 4782 565938 4866 566174
rect 5102 565938 44546 566174
rect 44782 565938 44866 566174
rect 45102 565938 84546 566174
rect 84782 565938 84866 566174
rect 85102 565938 124546 566174
rect 124782 565938 124866 566174
rect 125102 565938 164546 566174
rect 164782 565938 164866 566174
rect 165102 565938 204546 566174
rect 204782 565938 204866 566174
rect 205102 565938 244546 566174
rect 244782 565938 244866 566174
rect 245102 565938 284546 566174
rect 284782 565938 284866 566174
rect 285102 565938 324546 566174
rect 324782 565938 324866 566174
rect 325102 565938 364546 566174
rect 364782 565938 364866 566174
rect 365102 565938 404546 566174
rect 404782 565938 404866 566174
rect 405102 565938 444546 566174
rect 444782 565938 444866 566174
rect 445102 565938 484546 566174
rect 484782 565938 484866 566174
rect 485102 565938 524546 566174
rect 524782 565938 524866 566174
rect 525102 565938 564546 566174
rect 564782 565938 564866 566174
rect 565102 565938 587262 566174
rect 587498 565938 587582 566174
rect 587818 565938 588810 566174
rect -4886 565854 588810 565938
rect -4886 565618 -3894 565854
rect -3658 565618 -3574 565854
rect -3338 565618 4546 565854
rect 4782 565618 4866 565854
rect 5102 565618 44546 565854
rect 44782 565618 44866 565854
rect 45102 565618 84546 565854
rect 84782 565618 84866 565854
rect 85102 565618 124546 565854
rect 124782 565618 124866 565854
rect 125102 565618 164546 565854
rect 164782 565618 164866 565854
rect 165102 565618 204546 565854
rect 204782 565618 204866 565854
rect 205102 565618 244546 565854
rect 244782 565618 244866 565854
rect 245102 565618 284546 565854
rect 284782 565618 284866 565854
rect 285102 565618 324546 565854
rect 324782 565618 324866 565854
rect 325102 565618 364546 565854
rect 364782 565618 364866 565854
rect 365102 565618 404546 565854
rect 404782 565618 404866 565854
rect 405102 565618 444546 565854
rect 444782 565618 444866 565854
rect 445102 565618 484546 565854
rect 484782 565618 484866 565854
rect 485102 565618 524546 565854
rect 524782 565618 524866 565854
rect 525102 565618 564546 565854
rect 564782 565618 564866 565854
rect 565102 565618 587262 565854
rect 587498 565618 587582 565854
rect 587818 565618 588810 565854
rect -4886 565586 588810 565618
rect -2966 562454 586890 562486
rect -2966 562218 -1974 562454
rect -1738 562218 -1654 562454
rect -1418 562218 826 562454
rect 1062 562218 1146 562454
rect 1382 562218 40826 562454
rect 41062 562218 41146 562454
rect 41382 562218 80826 562454
rect 81062 562218 81146 562454
rect 81382 562218 120826 562454
rect 121062 562218 121146 562454
rect 121382 562218 160826 562454
rect 161062 562218 161146 562454
rect 161382 562218 200826 562454
rect 201062 562218 201146 562454
rect 201382 562218 240826 562454
rect 241062 562218 241146 562454
rect 241382 562218 280826 562454
rect 281062 562218 281146 562454
rect 281382 562218 320826 562454
rect 321062 562218 321146 562454
rect 321382 562218 360826 562454
rect 361062 562218 361146 562454
rect 361382 562218 400826 562454
rect 401062 562218 401146 562454
rect 401382 562218 440826 562454
rect 441062 562218 441146 562454
rect 441382 562218 480826 562454
rect 481062 562218 481146 562454
rect 481382 562218 520826 562454
rect 521062 562218 521146 562454
rect 521382 562218 560826 562454
rect 561062 562218 561146 562454
rect 561382 562218 585342 562454
rect 585578 562218 585662 562454
rect 585898 562218 586890 562454
rect -2966 562134 586890 562218
rect -2966 561898 -1974 562134
rect -1738 561898 -1654 562134
rect -1418 561898 826 562134
rect 1062 561898 1146 562134
rect 1382 561898 40826 562134
rect 41062 561898 41146 562134
rect 41382 561898 80826 562134
rect 81062 561898 81146 562134
rect 81382 561898 120826 562134
rect 121062 561898 121146 562134
rect 121382 561898 160826 562134
rect 161062 561898 161146 562134
rect 161382 561898 200826 562134
rect 201062 561898 201146 562134
rect 201382 561898 240826 562134
rect 241062 561898 241146 562134
rect 241382 561898 280826 562134
rect 281062 561898 281146 562134
rect 281382 561898 320826 562134
rect 321062 561898 321146 562134
rect 321382 561898 360826 562134
rect 361062 561898 361146 562134
rect 361382 561898 400826 562134
rect 401062 561898 401146 562134
rect 401382 561898 440826 562134
rect 441062 561898 441146 562134
rect 441382 561898 480826 562134
rect 481062 561898 481146 562134
rect 481382 561898 520826 562134
rect 521062 561898 521146 562134
rect 521382 561898 560826 562134
rect 561062 561898 561146 562134
rect 561382 561898 585342 562134
rect 585578 561898 585662 562134
rect 585898 561898 586890 562134
rect -2966 561866 586890 561898
rect -8726 553614 592650 553646
rect -8726 553378 -8694 553614
rect -8458 553378 -8374 553614
rect -8138 553378 31986 553614
rect 32222 553378 32306 553614
rect 32542 553378 71986 553614
rect 72222 553378 72306 553614
rect 72542 553378 111986 553614
rect 112222 553378 112306 553614
rect 112542 553378 151986 553614
rect 152222 553378 152306 553614
rect 152542 553378 191986 553614
rect 192222 553378 192306 553614
rect 192542 553378 231986 553614
rect 232222 553378 232306 553614
rect 232542 553378 271986 553614
rect 272222 553378 272306 553614
rect 272542 553378 311986 553614
rect 312222 553378 312306 553614
rect 312542 553378 351986 553614
rect 352222 553378 352306 553614
rect 352542 553378 391986 553614
rect 392222 553378 392306 553614
rect 392542 553378 431986 553614
rect 432222 553378 432306 553614
rect 432542 553378 471986 553614
rect 472222 553378 472306 553614
rect 472542 553378 511986 553614
rect 512222 553378 512306 553614
rect 512542 553378 551986 553614
rect 552222 553378 552306 553614
rect 552542 553378 592062 553614
rect 592298 553378 592382 553614
rect 592618 553378 592650 553614
rect -8726 553294 592650 553378
rect -8726 553058 -8694 553294
rect -8458 553058 -8374 553294
rect -8138 553058 31986 553294
rect 32222 553058 32306 553294
rect 32542 553058 71986 553294
rect 72222 553058 72306 553294
rect 72542 553058 111986 553294
rect 112222 553058 112306 553294
rect 112542 553058 151986 553294
rect 152222 553058 152306 553294
rect 152542 553058 191986 553294
rect 192222 553058 192306 553294
rect 192542 553058 231986 553294
rect 232222 553058 232306 553294
rect 232542 553058 271986 553294
rect 272222 553058 272306 553294
rect 272542 553058 311986 553294
rect 312222 553058 312306 553294
rect 312542 553058 351986 553294
rect 352222 553058 352306 553294
rect 352542 553058 391986 553294
rect 392222 553058 392306 553294
rect 392542 553058 431986 553294
rect 432222 553058 432306 553294
rect 432542 553058 471986 553294
rect 472222 553058 472306 553294
rect 472542 553058 511986 553294
rect 512222 553058 512306 553294
rect 512542 553058 551986 553294
rect 552222 553058 552306 553294
rect 552542 553058 592062 553294
rect 592298 553058 592382 553294
rect 592618 553058 592650 553294
rect -8726 553026 592650 553058
rect -6806 549894 590730 549926
rect -6806 549658 -6774 549894
rect -6538 549658 -6454 549894
rect -6218 549658 28266 549894
rect 28502 549658 28586 549894
rect 28822 549658 68266 549894
rect 68502 549658 68586 549894
rect 68822 549658 108266 549894
rect 108502 549658 108586 549894
rect 108822 549658 148266 549894
rect 148502 549658 148586 549894
rect 148822 549658 188266 549894
rect 188502 549658 188586 549894
rect 188822 549658 228266 549894
rect 228502 549658 228586 549894
rect 228822 549658 268266 549894
rect 268502 549658 268586 549894
rect 268822 549658 308266 549894
rect 308502 549658 308586 549894
rect 308822 549658 348266 549894
rect 348502 549658 348586 549894
rect 348822 549658 388266 549894
rect 388502 549658 388586 549894
rect 388822 549658 428266 549894
rect 428502 549658 428586 549894
rect 428822 549658 468266 549894
rect 468502 549658 468586 549894
rect 468822 549658 508266 549894
rect 508502 549658 508586 549894
rect 508822 549658 548266 549894
rect 548502 549658 548586 549894
rect 548822 549658 590142 549894
rect 590378 549658 590462 549894
rect 590698 549658 590730 549894
rect -6806 549574 590730 549658
rect -6806 549338 -6774 549574
rect -6538 549338 -6454 549574
rect -6218 549338 28266 549574
rect 28502 549338 28586 549574
rect 28822 549338 68266 549574
rect 68502 549338 68586 549574
rect 68822 549338 108266 549574
rect 108502 549338 108586 549574
rect 108822 549338 148266 549574
rect 148502 549338 148586 549574
rect 148822 549338 188266 549574
rect 188502 549338 188586 549574
rect 188822 549338 228266 549574
rect 228502 549338 228586 549574
rect 228822 549338 268266 549574
rect 268502 549338 268586 549574
rect 268822 549338 308266 549574
rect 308502 549338 308586 549574
rect 308822 549338 348266 549574
rect 348502 549338 348586 549574
rect 348822 549338 388266 549574
rect 388502 549338 388586 549574
rect 388822 549338 428266 549574
rect 428502 549338 428586 549574
rect 428822 549338 468266 549574
rect 468502 549338 468586 549574
rect 468822 549338 508266 549574
rect 508502 549338 508586 549574
rect 508822 549338 548266 549574
rect 548502 549338 548586 549574
rect 548822 549338 590142 549574
rect 590378 549338 590462 549574
rect 590698 549338 590730 549574
rect -6806 549306 590730 549338
rect -4886 546174 588810 546206
rect -4886 545938 -4854 546174
rect -4618 545938 -4534 546174
rect -4298 545938 24546 546174
rect 24782 545938 24866 546174
rect 25102 545938 64546 546174
rect 64782 545938 64866 546174
rect 65102 545938 104546 546174
rect 104782 545938 104866 546174
rect 105102 545938 144546 546174
rect 144782 545938 144866 546174
rect 145102 545938 184546 546174
rect 184782 545938 184866 546174
rect 185102 545938 224546 546174
rect 224782 545938 224866 546174
rect 225102 545938 264546 546174
rect 264782 545938 264866 546174
rect 265102 545938 304546 546174
rect 304782 545938 304866 546174
rect 305102 545938 344546 546174
rect 344782 545938 344866 546174
rect 345102 545938 384546 546174
rect 384782 545938 384866 546174
rect 385102 545938 424546 546174
rect 424782 545938 424866 546174
rect 425102 545938 464546 546174
rect 464782 545938 464866 546174
rect 465102 545938 504546 546174
rect 504782 545938 504866 546174
rect 505102 545938 544546 546174
rect 544782 545938 544866 546174
rect 545102 545938 588222 546174
rect 588458 545938 588542 546174
rect 588778 545938 588810 546174
rect -4886 545854 588810 545938
rect -4886 545618 -4854 545854
rect -4618 545618 -4534 545854
rect -4298 545618 24546 545854
rect 24782 545618 24866 545854
rect 25102 545618 64546 545854
rect 64782 545618 64866 545854
rect 65102 545618 104546 545854
rect 104782 545618 104866 545854
rect 105102 545618 144546 545854
rect 144782 545618 144866 545854
rect 145102 545618 184546 545854
rect 184782 545618 184866 545854
rect 185102 545618 224546 545854
rect 224782 545618 224866 545854
rect 225102 545618 264546 545854
rect 264782 545618 264866 545854
rect 265102 545618 304546 545854
rect 304782 545618 304866 545854
rect 305102 545618 344546 545854
rect 344782 545618 344866 545854
rect 345102 545618 384546 545854
rect 384782 545618 384866 545854
rect 385102 545618 424546 545854
rect 424782 545618 424866 545854
rect 425102 545618 464546 545854
rect 464782 545618 464866 545854
rect 465102 545618 504546 545854
rect 504782 545618 504866 545854
rect 505102 545618 544546 545854
rect 544782 545618 544866 545854
rect 545102 545618 588222 545854
rect 588458 545618 588542 545854
rect 588778 545618 588810 545854
rect -4886 545586 588810 545618
rect -2966 542454 586890 542486
rect -2966 542218 -2934 542454
rect -2698 542218 -2614 542454
rect -2378 542218 20826 542454
rect 21062 542218 21146 542454
rect 21382 542218 60826 542454
rect 61062 542218 61146 542454
rect 61382 542218 100826 542454
rect 101062 542218 101146 542454
rect 101382 542218 140826 542454
rect 141062 542218 141146 542454
rect 141382 542218 180826 542454
rect 181062 542218 181146 542454
rect 181382 542218 220826 542454
rect 221062 542218 221146 542454
rect 221382 542218 260826 542454
rect 261062 542218 261146 542454
rect 261382 542218 300826 542454
rect 301062 542218 301146 542454
rect 301382 542218 340826 542454
rect 341062 542218 341146 542454
rect 341382 542218 380826 542454
rect 381062 542218 381146 542454
rect 381382 542218 420826 542454
rect 421062 542218 421146 542454
rect 421382 542218 460826 542454
rect 461062 542218 461146 542454
rect 461382 542218 500826 542454
rect 501062 542218 501146 542454
rect 501382 542218 540826 542454
rect 541062 542218 541146 542454
rect 541382 542218 580826 542454
rect 581062 542218 581146 542454
rect 581382 542218 586302 542454
rect 586538 542218 586622 542454
rect 586858 542218 586890 542454
rect -2966 542134 586890 542218
rect -2966 541898 -2934 542134
rect -2698 541898 -2614 542134
rect -2378 541898 20826 542134
rect 21062 541898 21146 542134
rect 21382 541898 60826 542134
rect 61062 541898 61146 542134
rect 61382 541898 100826 542134
rect 101062 541898 101146 542134
rect 101382 541898 140826 542134
rect 141062 541898 141146 542134
rect 141382 541898 180826 542134
rect 181062 541898 181146 542134
rect 181382 541898 220826 542134
rect 221062 541898 221146 542134
rect 221382 541898 260826 542134
rect 261062 541898 261146 542134
rect 261382 541898 300826 542134
rect 301062 541898 301146 542134
rect 301382 541898 340826 542134
rect 341062 541898 341146 542134
rect 341382 541898 380826 542134
rect 381062 541898 381146 542134
rect 381382 541898 420826 542134
rect 421062 541898 421146 542134
rect 421382 541898 460826 542134
rect 461062 541898 461146 542134
rect 461382 541898 500826 542134
rect 501062 541898 501146 542134
rect 501382 541898 540826 542134
rect 541062 541898 541146 542134
rect 541382 541898 580826 542134
rect 581062 541898 581146 542134
rect 581382 541898 586302 542134
rect 586538 541898 586622 542134
rect 586858 541898 586890 542134
rect -2966 541866 586890 541898
rect -8726 533614 592650 533646
rect -8726 533378 -7734 533614
rect -7498 533378 -7414 533614
rect -7178 533378 11986 533614
rect 12222 533378 12306 533614
rect 12542 533378 51986 533614
rect 52222 533378 52306 533614
rect 52542 533378 91986 533614
rect 92222 533378 92306 533614
rect 92542 533378 131986 533614
rect 132222 533378 132306 533614
rect 132542 533378 171986 533614
rect 172222 533378 172306 533614
rect 172542 533378 211986 533614
rect 212222 533378 212306 533614
rect 212542 533378 251986 533614
rect 252222 533378 252306 533614
rect 252542 533378 291986 533614
rect 292222 533378 292306 533614
rect 292542 533378 331986 533614
rect 332222 533378 332306 533614
rect 332542 533378 371986 533614
rect 372222 533378 372306 533614
rect 372542 533378 411986 533614
rect 412222 533378 412306 533614
rect 412542 533378 451986 533614
rect 452222 533378 452306 533614
rect 452542 533378 491986 533614
rect 492222 533378 492306 533614
rect 492542 533378 531986 533614
rect 532222 533378 532306 533614
rect 532542 533378 571986 533614
rect 572222 533378 572306 533614
rect 572542 533378 591102 533614
rect 591338 533378 591422 533614
rect 591658 533378 592650 533614
rect -8726 533294 592650 533378
rect -8726 533058 -7734 533294
rect -7498 533058 -7414 533294
rect -7178 533058 11986 533294
rect 12222 533058 12306 533294
rect 12542 533058 51986 533294
rect 52222 533058 52306 533294
rect 52542 533058 91986 533294
rect 92222 533058 92306 533294
rect 92542 533058 131986 533294
rect 132222 533058 132306 533294
rect 132542 533058 171986 533294
rect 172222 533058 172306 533294
rect 172542 533058 211986 533294
rect 212222 533058 212306 533294
rect 212542 533058 251986 533294
rect 252222 533058 252306 533294
rect 252542 533058 291986 533294
rect 292222 533058 292306 533294
rect 292542 533058 331986 533294
rect 332222 533058 332306 533294
rect 332542 533058 371986 533294
rect 372222 533058 372306 533294
rect 372542 533058 411986 533294
rect 412222 533058 412306 533294
rect 412542 533058 451986 533294
rect 452222 533058 452306 533294
rect 452542 533058 491986 533294
rect 492222 533058 492306 533294
rect 492542 533058 531986 533294
rect 532222 533058 532306 533294
rect 532542 533058 571986 533294
rect 572222 533058 572306 533294
rect 572542 533058 591102 533294
rect 591338 533058 591422 533294
rect 591658 533058 592650 533294
rect -8726 533026 592650 533058
rect -6806 529894 590730 529926
rect -6806 529658 -5814 529894
rect -5578 529658 -5494 529894
rect -5258 529658 8266 529894
rect 8502 529658 8586 529894
rect 8822 529658 48266 529894
rect 48502 529658 48586 529894
rect 48822 529658 88266 529894
rect 88502 529658 88586 529894
rect 88822 529658 128266 529894
rect 128502 529658 128586 529894
rect 128822 529658 168266 529894
rect 168502 529658 168586 529894
rect 168822 529658 208266 529894
rect 208502 529658 208586 529894
rect 208822 529658 248266 529894
rect 248502 529658 248586 529894
rect 248822 529658 288266 529894
rect 288502 529658 288586 529894
rect 288822 529658 328266 529894
rect 328502 529658 328586 529894
rect 328822 529658 368266 529894
rect 368502 529658 368586 529894
rect 368822 529658 408266 529894
rect 408502 529658 408586 529894
rect 408822 529658 448266 529894
rect 448502 529658 448586 529894
rect 448822 529658 488266 529894
rect 488502 529658 488586 529894
rect 488822 529658 528266 529894
rect 528502 529658 528586 529894
rect 528822 529658 568266 529894
rect 568502 529658 568586 529894
rect 568822 529658 589182 529894
rect 589418 529658 589502 529894
rect 589738 529658 590730 529894
rect -6806 529574 590730 529658
rect -6806 529338 -5814 529574
rect -5578 529338 -5494 529574
rect -5258 529338 8266 529574
rect 8502 529338 8586 529574
rect 8822 529338 48266 529574
rect 48502 529338 48586 529574
rect 48822 529338 88266 529574
rect 88502 529338 88586 529574
rect 88822 529338 128266 529574
rect 128502 529338 128586 529574
rect 128822 529338 168266 529574
rect 168502 529338 168586 529574
rect 168822 529338 208266 529574
rect 208502 529338 208586 529574
rect 208822 529338 248266 529574
rect 248502 529338 248586 529574
rect 248822 529338 288266 529574
rect 288502 529338 288586 529574
rect 288822 529338 328266 529574
rect 328502 529338 328586 529574
rect 328822 529338 368266 529574
rect 368502 529338 368586 529574
rect 368822 529338 408266 529574
rect 408502 529338 408586 529574
rect 408822 529338 448266 529574
rect 448502 529338 448586 529574
rect 448822 529338 488266 529574
rect 488502 529338 488586 529574
rect 488822 529338 528266 529574
rect 528502 529338 528586 529574
rect 528822 529338 568266 529574
rect 568502 529338 568586 529574
rect 568822 529338 589182 529574
rect 589418 529338 589502 529574
rect 589738 529338 590730 529574
rect -6806 529306 590730 529338
rect -4886 526174 588810 526206
rect -4886 525938 -3894 526174
rect -3658 525938 -3574 526174
rect -3338 525938 4546 526174
rect 4782 525938 4866 526174
rect 5102 525938 44546 526174
rect 44782 525938 44866 526174
rect 45102 525938 84546 526174
rect 84782 525938 84866 526174
rect 85102 525938 124546 526174
rect 124782 525938 124866 526174
rect 125102 525938 164546 526174
rect 164782 525938 164866 526174
rect 165102 525938 204546 526174
rect 204782 525938 204866 526174
rect 205102 525938 244546 526174
rect 244782 525938 244866 526174
rect 245102 525938 284546 526174
rect 284782 525938 284866 526174
rect 285102 525938 324546 526174
rect 324782 525938 324866 526174
rect 325102 525938 364546 526174
rect 364782 525938 364866 526174
rect 365102 525938 404546 526174
rect 404782 525938 404866 526174
rect 405102 525938 444546 526174
rect 444782 525938 444866 526174
rect 445102 525938 484546 526174
rect 484782 525938 484866 526174
rect 485102 525938 524546 526174
rect 524782 525938 524866 526174
rect 525102 525938 564546 526174
rect 564782 525938 564866 526174
rect 565102 525938 587262 526174
rect 587498 525938 587582 526174
rect 587818 525938 588810 526174
rect -4886 525854 588810 525938
rect -4886 525618 -3894 525854
rect -3658 525618 -3574 525854
rect -3338 525618 4546 525854
rect 4782 525618 4866 525854
rect 5102 525618 44546 525854
rect 44782 525618 44866 525854
rect 45102 525618 84546 525854
rect 84782 525618 84866 525854
rect 85102 525618 124546 525854
rect 124782 525618 124866 525854
rect 125102 525618 164546 525854
rect 164782 525618 164866 525854
rect 165102 525618 204546 525854
rect 204782 525618 204866 525854
rect 205102 525618 244546 525854
rect 244782 525618 244866 525854
rect 245102 525618 284546 525854
rect 284782 525618 284866 525854
rect 285102 525618 324546 525854
rect 324782 525618 324866 525854
rect 325102 525618 364546 525854
rect 364782 525618 364866 525854
rect 365102 525618 404546 525854
rect 404782 525618 404866 525854
rect 405102 525618 444546 525854
rect 444782 525618 444866 525854
rect 445102 525618 484546 525854
rect 484782 525618 484866 525854
rect 485102 525618 524546 525854
rect 524782 525618 524866 525854
rect 525102 525618 564546 525854
rect 564782 525618 564866 525854
rect 565102 525618 587262 525854
rect 587498 525618 587582 525854
rect 587818 525618 588810 525854
rect -4886 525586 588810 525618
rect -2966 522454 586890 522486
rect -2966 522218 -1974 522454
rect -1738 522218 -1654 522454
rect -1418 522218 826 522454
rect 1062 522218 1146 522454
rect 1382 522218 40826 522454
rect 41062 522218 41146 522454
rect 41382 522218 80826 522454
rect 81062 522218 81146 522454
rect 81382 522218 120826 522454
rect 121062 522218 121146 522454
rect 121382 522218 160826 522454
rect 161062 522218 161146 522454
rect 161382 522218 200826 522454
rect 201062 522218 201146 522454
rect 201382 522218 240826 522454
rect 241062 522218 241146 522454
rect 241382 522218 280826 522454
rect 281062 522218 281146 522454
rect 281382 522218 320826 522454
rect 321062 522218 321146 522454
rect 321382 522218 360826 522454
rect 361062 522218 361146 522454
rect 361382 522218 400826 522454
rect 401062 522218 401146 522454
rect 401382 522218 440826 522454
rect 441062 522218 441146 522454
rect 441382 522218 480826 522454
rect 481062 522218 481146 522454
rect 481382 522218 520826 522454
rect 521062 522218 521146 522454
rect 521382 522218 560826 522454
rect 561062 522218 561146 522454
rect 561382 522218 585342 522454
rect 585578 522218 585662 522454
rect 585898 522218 586890 522454
rect -2966 522134 586890 522218
rect -2966 521898 -1974 522134
rect -1738 521898 -1654 522134
rect -1418 521898 826 522134
rect 1062 521898 1146 522134
rect 1382 521898 40826 522134
rect 41062 521898 41146 522134
rect 41382 521898 80826 522134
rect 81062 521898 81146 522134
rect 81382 521898 120826 522134
rect 121062 521898 121146 522134
rect 121382 521898 160826 522134
rect 161062 521898 161146 522134
rect 161382 521898 200826 522134
rect 201062 521898 201146 522134
rect 201382 521898 240826 522134
rect 241062 521898 241146 522134
rect 241382 521898 280826 522134
rect 281062 521898 281146 522134
rect 281382 521898 320826 522134
rect 321062 521898 321146 522134
rect 321382 521898 360826 522134
rect 361062 521898 361146 522134
rect 361382 521898 400826 522134
rect 401062 521898 401146 522134
rect 401382 521898 440826 522134
rect 441062 521898 441146 522134
rect 441382 521898 480826 522134
rect 481062 521898 481146 522134
rect 481382 521898 520826 522134
rect 521062 521898 521146 522134
rect 521382 521898 560826 522134
rect 561062 521898 561146 522134
rect 561382 521898 585342 522134
rect 585578 521898 585662 522134
rect 585898 521898 586890 522134
rect -2966 521866 586890 521898
rect -8726 513614 592650 513646
rect -8726 513378 -8694 513614
rect -8458 513378 -8374 513614
rect -8138 513378 31986 513614
rect 32222 513378 32306 513614
rect 32542 513378 71986 513614
rect 72222 513378 72306 513614
rect 72542 513378 111986 513614
rect 112222 513378 112306 513614
rect 112542 513378 151986 513614
rect 152222 513378 152306 513614
rect 152542 513378 191986 513614
rect 192222 513378 192306 513614
rect 192542 513378 231986 513614
rect 232222 513378 232306 513614
rect 232542 513378 271986 513614
rect 272222 513378 272306 513614
rect 272542 513378 311986 513614
rect 312222 513378 312306 513614
rect 312542 513378 351986 513614
rect 352222 513378 352306 513614
rect 352542 513378 391986 513614
rect 392222 513378 392306 513614
rect 392542 513378 431986 513614
rect 432222 513378 432306 513614
rect 432542 513378 471986 513614
rect 472222 513378 472306 513614
rect 472542 513378 511986 513614
rect 512222 513378 512306 513614
rect 512542 513378 551986 513614
rect 552222 513378 552306 513614
rect 552542 513378 592062 513614
rect 592298 513378 592382 513614
rect 592618 513378 592650 513614
rect -8726 513294 592650 513378
rect -8726 513058 -8694 513294
rect -8458 513058 -8374 513294
rect -8138 513058 31986 513294
rect 32222 513058 32306 513294
rect 32542 513058 71986 513294
rect 72222 513058 72306 513294
rect 72542 513058 111986 513294
rect 112222 513058 112306 513294
rect 112542 513058 151986 513294
rect 152222 513058 152306 513294
rect 152542 513058 191986 513294
rect 192222 513058 192306 513294
rect 192542 513058 231986 513294
rect 232222 513058 232306 513294
rect 232542 513058 271986 513294
rect 272222 513058 272306 513294
rect 272542 513058 311986 513294
rect 312222 513058 312306 513294
rect 312542 513058 351986 513294
rect 352222 513058 352306 513294
rect 352542 513058 391986 513294
rect 392222 513058 392306 513294
rect 392542 513058 431986 513294
rect 432222 513058 432306 513294
rect 432542 513058 471986 513294
rect 472222 513058 472306 513294
rect 472542 513058 511986 513294
rect 512222 513058 512306 513294
rect 512542 513058 551986 513294
rect 552222 513058 552306 513294
rect 552542 513058 592062 513294
rect 592298 513058 592382 513294
rect 592618 513058 592650 513294
rect -8726 513026 592650 513058
rect -6806 509894 590730 509926
rect -6806 509658 -6774 509894
rect -6538 509658 -6454 509894
rect -6218 509658 28266 509894
rect 28502 509658 28586 509894
rect 28822 509658 68266 509894
rect 68502 509658 68586 509894
rect 68822 509658 108266 509894
rect 108502 509658 108586 509894
rect 108822 509658 148266 509894
rect 148502 509658 148586 509894
rect 148822 509658 188266 509894
rect 188502 509658 188586 509894
rect 188822 509658 228266 509894
rect 228502 509658 228586 509894
rect 228822 509658 268266 509894
rect 268502 509658 268586 509894
rect 268822 509658 308266 509894
rect 308502 509658 308586 509894
rect 308822 509658 348266 509894
rect 348502 509658 348586 509894
rect 348822 509658 388266 509894
rect 388502 509658 388586 509894
rect 388822 509658 428266 509894
rect 428502 509658 428586 509894
rect 428822 509658 468266 509894
rect 468502 509658 468586 509894
rect 468822 509658 508266 509894
rect 508502 509658 508586 509894
rect 508822 509658 548266 509894
rect 548502 509658 548586 509894
rect 548822 509658 590142 509894
rect 590378 509658 590462 509894
rect 590698 509658 590730 509894
rect -6806 509574 590730 509658
rect -6806 509338 -6774 509574
rect -6538 509338 -6454 509574
rect -6218 509338 28266 509574
rect 28502 509338 28586 509574
rect 28822 509338 68266 509574
rect 68502 509338 68586 509574
rect 68822 509338 108266 509574
rect 108502 509338 108586 509574
rect 108822 509338 148266 509574
rect 148502 509338 148586 509574
rect 148822 509338 188266 509574
rect 188502 509338 188586 509574
rect 188822 509338 228266 509574
rect 228502 509338 228586 509574
rect 228822 509338 268266 509574
rect 268502 509338 268586 509574
rect 268822 509338 308266 509574
rect 308502 509338 308586 509574
rect 308822 509338 348266 509574
rect 348502 509338 348586 509574
rect 348822 509338 388266 509574
rect 388502 509338 388586 509574
rect 388822 509338 428266 509574
rect 428502 509338 428586 509574
rect 428822 509338 468266 509574
rect 468502 509338 468586 509574
rect 468822 509338 508266 509574
rect 508502 509338 508586 509574
rect 508822 509338 548266 509574
rect 548502 509338 548586 509574
rect 548822 509338 590142 509574
rect 590378 509338 590462 509574
rect 590698 509338 590730 509574
rect -6806 509306 590730 509338
rect -4886 506174 588810 506206
rect -4886 505938 -4854 506174
rect -4618 505938 -4534 506174
rect -4298 505938 24546 506174
rect 24782 505938 24866 506174
rect 25102 505938 64546 506174
rect 64782 505938 64866 506174
rect 65102 505938 104546 506174
rect 104782 505938 104866 506174
rect 105102 505938 144546 506174
rect 144782 505938 144866 506174
rect 145102 505938 184546 506174
rect 184782 505938 184866 506174
rect 185102 505938 224546 506174
rect 224782 505938 224866 506174
rect 225102 505938 264546 506174
rect 264782 505938 264866 506174
rect 265102 505938 304546 506174
rect 304782 505938 304866 506174
rect 305102 505938 344546 506174
rect 344782 505938 344866 506174
rect 345102 505938 384546 506174
rect 384782 505938 384866 506174
rect 385102 505938 424546 506174
rect 424782 505938 424866 506174
rect 425102 505938 464546 506174
rect 464782 505938 464866 506174
rect 465102 505938 504546 506174
rect 504782 505938 504866 506174
rect 505102 505938 544546 506174
rect 544782 505938 544866 506174
rect 545102 505938 588222 506174
rect 588458 505938 588542 506174
rect 588778 505938 588810 506174
rect -4886 505854 588810 505938
rect -4886 505618 -4854 505854
rect -4618 505618 -4534 505854
rect -4298 505618 24546 505854
rect 24782 505618 24866 505854
rect 25102 505618 64546 505854
rect 64782 505618 64866 505854
rect 65102 505618 104546 505854
rect 104782 505618 104866 505854
rect 105102 505618 144546 505854
rect 144782 505618 144866 505854
rect 145102 505618 184546 505854
rect 184782 505618 184866 505854
rect 185102 505618 224546 505854
rect 224782 505618 224866 505854
rect 225102 505618 264546 505854
rect 264782 505618 264866 505854
rect 265102 505618 304546 505854
rect 304782 505618 304866 505854
rect 305102 505618 344546 505854
rect 344782 505618 344866 505854
rect 345102 505618 384546 505854
rect 384782 505618 384866 505854
rect 385102 505618 424546 505854
rect 424782 505618 424866 505854
rect 425102 505618 464546 505854
rect 464782 505618 464866 505854
rect 465102 505618 504546 505854
rect 504782 505618 504866 505854
rect 505102 505618 544546 505854
rect 544782 505618 544866 505854
rect 545102 505618 588222 505854
rect 588458 505618 588542 505854
rect 588778 505618 588810 505854
rect -4886 505586 588810 505618
rect -2966 502454 586890 502486
rect -2966 502218 -2934 502454
rect -2698 502218 -2614 502454
rect -2378 502218 20826 502454
rect 21062 502218 21146 502454
rect 21382 502218 60826 502454
rect 61062 502218 61146 502454
rect 61382 502218 100826 502454
rect 101062 502218 101146 502454
rect 101382 502218 140826 502454
rect 141062 502218 141146 502454
rect 141382 502218 180826 502454
rect 181062 502218 181146 502454
rect 181382 502218 220826 502454
rect 221062 502218 221146 502454
rect 221382 502218 260826 502454
rect 261062 502218 261146 502454
rect 261382 502218 300826 502454
rect 301062 502218 301146 502454
rect 301382 502218 340826 502454
rect 341062 502218 341146 502454
rect 341382 502218 380826 502454
rect 381062 502218 381146 502454
rect 381382 502218 420826 502454
rect 421062 502218 421146 502454
rect 421382 502218 460826 502454
rect 461062 502218 461146 502454
rect 461382 502218 500826 502454
rect 501062 502218 501146 502454
rect 501382 502218 540826 502454
rect 541062 502218 541146 502454
rect 541382 502218 580826 502454
rect 581062 502218 581146 502454
rect 581382 502218 586302 502454
rect 586538 502218 586622 502454
rect 586858 502218 586890 502454
rect -2966 502134 586890 502218
rect -2966 501898 -2934 502134
rect -2698 501898 -2614 502134
rect -2378 501898 20826 502134
rect 21062 501898 21146 502134
rect 21382 501898 60826 502134
rect 61062 501898 61146 502134
rect 61382 501898 100826 502134
rect 101062 501898 101146 502134
rect 101382 501898 140826 502134
rect 141062 501898 141146 502134
rect 141382 501898 180826 502134
rect 181062 501898 181146 502134
rect 181382 501898 220826 502134
rect 221062 501898 221146 502134
rect 221382 501898 260826 502134
rect 261062 501898 261146 502134
rect 261382 501898 300826 502134
rect 301062 501898 301146 502134
rect 301382 501898 340826 502134
rect 341062 501898 341146 502134
rect 341382 501898 380826 502134
rect 381062 501898 381146 502134
rect 381382 501898 420826 502134
rect 421062 501898 421146 502134
rect 421382 501898 460826 502134
rect 461062 501898 461146 502134
rect 461382 501898 500826 502134
rect 501062 501898 501146 502134
rect 501382 501898 540826 502134
rect 541062 501898 541146 502134
rect 541382 501898 580826 502134
rect 581062 501898 581146 502134
rect 581382 501898 586302 502134
rect 586538 501898 586622 502134
rect 586858 501898 586890 502134
rect -2966 501866 586890 501898
rect -8726 493614 592650 493646
rect -8726 493378 -7734 493614
rect -7498 493378 -7414 493614
rect -7178 493378 11986 493614
rect 12222 493378 12306 493614
rect 12542 493378 51986 493614
rect 52222 493378 52306 493614
rect 52542 493378 91986 493614
rect 92222 493378 92306 493614
rect 92542 493378 131986 493614
rect 132222 493378 132306 493614
rect 132542 493378 171986 493614
rect 172222 493378 172306 493614
rect 172542 493378 211986 493614
rect 212222 493378 212306 493614
rect 212542 493378 251986 493614
rect 252222 493378 252306 493614
rect 252542 493378 291986 493614
rect 292222 493378 292306 493614
rect 292542 493378 331986 493614
rect 332222 493378 332306 493614
rect 332542 493378 371986 493614
rect 372222 493378 372306 493614
rect 372542 493378 411986 493614
rect 412222 493378 412306 493614
rect 412542 493378 451986 493614
rect 452222 493378 452306 493614
rect 452542 493378 491986 493614
rect 492222 493378 492306 493614
rect 492542 493378 531986 493614
rect 532222 493378 532306 493614
rect 532542 493378 571986 493614
rect 572222 493378 572306 493614
rect 572542 493378 591102 493614
rect 591338 493378 591422 493614
rect 591658 493378 592650 493614
rect -8726 493294 592650 493378
rect -8726 493058 -7734 493294
rect -7498 493058 -7414 493294
rect -7178 493058 11986 493294
rect 12222 493058 12306 493294
rect 12542 493058 51986 493294
rect 52222 493058 52306 493294
rect 52542 493058 91986 493294
rect 92222 493058 92306 493294
rect 92542 493058 131986 493294
rect 132222 493058 132306 493294
rect 132542 493058 171986 493294
rect 172222 493058 172306 493294
rect 172542 493058 211986 493294
rect 212222 493058 212306 493294
rect 212542 493058 251986 493294
rect 252222 493058 252306 493294
rect 252542 493058 291986 493294
rect 292222 493058 292306 493294
rect 292542 493058 331986 493294
rect 332222 493058 332306 493294
rect 332542 493058 371986 493294
rect 372222 493058 372306 493294
rect 372542 493058 411986 493294
rect 412222 493058 412306 493294
rect 412542 493058 451986 493294
rect 452222 493058 452306 493294
rect 452542 493058 491986 493294
rect 492222 493058 492306 493294
rect 492542 493058 531986 493294
rect 532222 493058 532306 493294
rect 532542 493058 571986 493294
rect 572222 493058 572306 493294
rect 572542 493058 591102 493294
rect 591338 493058 591422 493294
rect 591658 493058 592650 493294
rect -8726 493026 592650 493058
rect -6806 489894 590730 489926
rect -6806 489658 -5814 489894
rect -5578 489658 -5494 489894
rect -5258 489658 8266 489894
rect 8502 489658 8586 489894
rect 8822 489658 48266 489894
rect 48502 489658 48586 489894
rect 48822 489658 88266 489894
rect 88502 489658 88586 489894
rect 88822 489658 128266 489894
rect 128502 489658 128586 489894
rect 128822 489658 168266 489894
rect 168502 489658 168586 489894
rect 168822 489658 208266 489894
rect 208502 489658 208586 489894
rect 208822 489658 248266 489894
rect 248502 489658 248586 489894
rect 248822 489658 288266 489894
rect 288502 489658 288586 489894
rect 288822 489658 328266 489894
rect 328502 489658 328586 489894
rect 328822 489658 368266 489894
rect 368502 489658 368586 489894
rect 368822 489658 408266 489894
rect 408502 489658 408586 489894
rect 408822 489658 448266 489894
rect 448502 489658 448586 489894
rect 448822 489658 488266 489894
rect 488502 489658 488586 489894
rect 488822 489658 528266 489894
rect 528502 489658 528586 489894
rect 528822 489658 568266 489894
rect 568502 489658 568586 489894
rect 568822 489658 589182 489894
rect 589418 489658 589502 489894
rect 589738 489658 590730 489894
rect -6806 489574 590730 489658
rect -6806 489338 -5814 489574
rect -5578 489338 -5494 489574
rect -5258 489338 8266 489574
rect 8502 489338 8586 489574
rect 8822 489338 48266 489574
rect 48502 489338 48586 489574
rect 48822 489338 88266 489574
rect 88502 489338 88586 489574
rect 88822 489338 128266 489574
rect 128502 489338 128586 489574
rect 128822 489338 168266 489574
rect 168502 489338 168586 489574
rect 168822 489338 208266 489574
rect 208502 489338 208586 489574
rect 208822 489338 248266 489574
rect 248502 489338 248586 489574
rect 248822 489338 288266 489574
rect 288502 489338 288586 489574
rect 288822 489338 328266 489574
rect 328502 489338 328586 489574
rect 328822 489338 368266 489574
rect 368502 489338 368586 489574
rect 368822 489338 408266 489574
rect 408502 489338 408586 489574
rect 408822 489338 448266 489574
rect 448502 489338 448586 489574
rect 448822 489338 488266 489574
rect 488502 489338 488586 489574
rect 488822 489338 528266 489574
rect 528502 489338 528586 489574
rect 528822 489338 568266 489574
rect 568502 489338 568586 489574
rect 568822 489338 589182 489574
rect 589418 489338 589502 489574
rect 589738 489338 590730 489574
rect -6806 489306 590730 489338
rect -4886 486174 588810 486206
rect -4886 485938 -3894 486174
rect -3658 485938 -3574 486174
rect -3338 485938 4546 486174
rect 4782 485938 4866 486174
rect 5102 485938 44546 486174
rect 44782 485938 44866 486174
rect 45102 485938 84546 486174
rect 84782 485938 84866 486174
rect 85102 485938 124546 486174
rect 124782 485938 124866 486174
rect 125102 485938 164546 486174
rect 164782 485938 164866 486174
rect 165102 485938 204546 486174
rect 204782 485938 204866 486174
rect 205102 485938 244546 486174
rect 244782 485938 244866 486174
rect 245102 485938 284546 486174
rect 284782 485938 284866 486174
rect 285102 485938 324546 486174
rect 324782 485938 324866 486174
rect 325102 485938 364546 486174
rect 364782 485938 364866 486174
rect 365102 485938 404546 486174
rect 404782 485938 404866 486174
rect 405102 485938 444546 486174
rect 444782 485938 444866 486174
rect 445102 485938 484546 486174
rect 484782 485938 484866 486174
rect 485102 485938 524546 486174
rect 524782 485938 524866 486174
rect 525102 485938 564546 486174
rect 564782 485938 564866 486174
rect 565102 485938 587262 486174
rect 587498 485938 587582 486174
rect 587818 485938 588810 486174
rect -4886 485854 588810 485938
rect -4886 485618 -3894 485854
rect -3658 485618 -3574 485854
rect -3338 485618 4546 485854
rect 4782 485618 4866 485854
rect 5102 485618 44546 485854
rect 44782 485618 44866 485854
rect 45102 485618 84546 485854
rect 84782 485618 84866 485854
rect 85102 485618 124546 485854
rect 124782 485618 124866 485854
rect 125102 485618 164546 485854
rect 164782 485618 164866 485854
rect 165102 485618 204546 485854
rect 204782 485618 204866 485854
rect 205102 485618 244546 485854
rect 244782 485618 244866 485854
rect 245102 485618 284546 485854
rect 284782 485618 284866 485854
rect 285102 485618 324546 485854
rect 324782 485618 324866 485854
rect 325102 485618 364546 485854
rect 364782 485618 364866 485854
rect 365102 485618 404546 485854
rect 404782 485618 404866 485854
rect 405102 485618 444546 485854
rect 444782 485618 444866 485854
rect 445102 485618 484546 485854
rect 484782 485618 484866 485854
rect 485102 485618 524546 485854
rect 524782 485618 524866 485854
rect 525102 485618 564546 485854
rect 564782 485618 564866 485854
rect 565102 485618 587262 485854
rect 587498 485618 587582 485854
rect 587818 485618 588810 485854
rect -4886 485586 588810 485618
rect -2966 482454 586890 482486
rect -2966 482218 -1974 482454
rect -1738 482218 -1654 482454
rect -1418 482218 826 482454
rect 1062 482218 1146 482454
rect 1382 482218 40826 482454
rect 41062 482218 41146 482454
rect 41382 482218 80826 482454
rect 81062 482218 81146 482454
rect 81382 482218 120826 482454
rect 121062 482218 121146 482454
rect 121382 482218 160826 482454
rect 161062 482218 161146 482454
rect 161382 482218 200826 482454
rect 201062 482218 201146 482454
rect 201382 482218 240826 482454
rect 241062 482218 241146 482454
rect 241382 482218 280826 482454
rect 281062 482218 281146 482454
rect 281382 482218 320826 482454
rect 321062 482218 321146 482454
rect 321382 482218 360826 482454
rect 361062 482218 361146 482454
rect 361382 482218 400826 482454
rect 401062 482218 401146 482454
rect 401382 482218 440826 482454
rect 441062 482218 441146 482454
rect 441382 482218 480826 482454
rect 481062 482218 481146 482454
rect 481382 482218 520826 482454
rect 521062 482218 521146 482454
rect 521382 482218 560826 482454
rect 561062 482218 561146 482454
rect 561382 482218 585342 482454
rect 585578 482218 585662 482454
rect 585898 482218 586890 482454
rect -2966 482134 586890 482218
rect -2966 481898 -1974 482134
rect -1738 481898 -1654 482134
rect -1418 481898 826 482134
rect 1062 481898 1146 482134
rect 1382 481898 40826 482134
rect 41062 481898 41146 482134
rect 41382 481898 80826 482134
rect 81062 481898 81146 482134
rect 81382 481898 120826 482134
rect 121062 481898 121146 482134
rect 121382 481898 160826 482134
rect 161062 481898 161146 482134
rect 161382 481898 200826 482134
rect 201062 481898 201146 482134
rect 201382 481898 240826 482134
rect 241062 481898 241146 482134
rect 241382 481898 280826 482134
rect 281062 481898 281146 482134
rect 281382 481898 320826 482134
rect 321062 481898 321146 482134
rect 321382 481898 360826 482134
rect 361062 481898 361146 482134
rect 361382 481898 400826 482134
rect 401062 481898 401146 482134
rect 401382 481898 440826 482134
rect 441062 481898 441146 482134
rect 441382 481898 480826 482134
rect 481062 481898 481146 482134
rect 481382 481898 520826 482134
rect 521062 481898 521146 482134
rect 521382 481898 560826 482134
rect 561062 481898 561146 482134
rect 561382 481898 585342 482134
rect 585578 481898 585662 482134
rect 585898 481898 586890 482134
rect -2966 481866 586890 481898
rect -8726 473614 592650 473646
rect -8726 473378 -8694 473614
rect -8458 473378 -8374 473614
rect -8138 473378 31986 473614
rect 32222 473378 32306 473614
rect 32542 473378 71986 473614
rect 72222 473378 72306 473614
rect 72542 473378 111986 473614
rect 112222 473378 112306 473614
rect 112542 473378 151986 473614
rect 152222 473378 152306 473614
rect 152542 473378 191986 473614
rect 192222 473378 192306 473614
rect 192542 473378 231986 473614
rect 232222 473378 232306 473614
rect 232542 473378 271986 473614
rect 272222 473378 272306 473614
rect 272542 473378 311986 473614
rect 312222 473378 312306 473614
rect 312542 473378 351986 473614
rect 352222 473378 352306 473614
rect 352542 473378 391986 473614
rect 392222 473378 392306 473614
rect 392542 473378 431986 473614
rect 432222 473378 432306 473614
rect 432542 473378 471986 473614
rect 472222 473378 472306 473614
rect 472542 473378 511986 473614
rect 512222 473378 512306 473614
rect 512542 473378 551986 473614
rect 552222 473378 552306 473614
rect 552542 473378 592062 473614
rect 592298 473378 592382 473614
rect 592618 473378 592650 473614
rect -8726 473294 592650 473378
rect -8726 473058 -8694 473294
rect -8458 473058 -8374 473294
rect -8138 473058 31986 473294
rect 32222 473058 32306 473294
rect 32542 473058 71986 473294
rect 72222 473058 72306 473294
rect 72542 473058 111986 473294
rect 112222 473058 112306 473294
rect 112542 473058 151986 473294
rect 152222 473058 152306 473294
rect 152542 473058 191986 473294
rect 192222 473058 192306 473294
rect 192542 473058 231986 473294
rect 232222 473058 232306 473294
rect 232542 473058 271986 473294
rect 272222 473058 272306 473294
rect 272542 473058 311986 473294
rect 312222 473058 312306 473294
rect 312542 473058 351986 473294
rect 352222 473058 352306 473294
rect 352542 473058 391986 473294
rect 392222 473058 392306 473294
rect 392542 473058 431986 473294
rect 432222 473058 432306 473294
rect 432542 473058 471986 473294
rect 472222 473058 472306 473294
rect 472542 473058 511986 473294
rect 512222 473058 512306 473294
rect 512542 473058 551986 473294
rect 552222 473058 552306 473294
rect 552542 473058 592062 473294
rect 592298 473058 592382 473294
rect 592618 473058 592650 473294
rect -8726 473026 592650 473058
rect -6806 469894 590730 469926
rect -6806 469658 -6774 469894
rect -6538 469658 -6454 469894
rect -6218 469658 28266 469894
rect 28502 469658 28586 469894
rect 28822 469658 68266 469894
rect 68502 469658 68586 469894
rect 68822 469658 108266 469894
rect 108502 469658 108586 469894
rect 108822 469658 148266 469894
rect 148502 469658 148586 469894
rect 148822 469658 188266 469894
rect 188502 469658 188586 469894
rect 188822 469658 228266 469894
rect 228502 469658 228586 469894
rect 228822 469658 268266 469894
rect 268502 469658 268586 469894
rect 268822 469658 308266 469894
rect 308502 469658 308586 469894
rect 308822 469658 348266 469894
rect 348502 469658 348586 469894
rect 348822 469658 388266 469894
rect 388502 469658 388586 469894
rect 388822 469658 428266 469894
rect 428502 469658 428586 469894
rect 428822 469658 468266 469894
rect 468502 469658 468586 469894
rect 468822 469658 508266 469894
rect 508502 469658 508586 469894
rect 508822 469658 548266 469894
rect 548502 469658 548586 469894
rect 548822 469658 590142 469894
rect 590378 469658 590462 469894
rect 590698 469658 590730 469894
rect -6806 469574 590730 469658
rect -6806 469338 -6774 469574
rect -6538 469338 -6454 469574
rect -6218 469338 28266 469574
rect 28502 469338 28586 469574
rect 28822 469338 68266 469574
rect 68502 469338 68586 469574
rect 68822 469338 108266 469574
rect 108502 469338 108586 469574
rect 108822 469338 148266 469574
rect 148502 469338 148586 469574
rect 148822 469338 188266 469574
rect 188502 469338 188586 469574
rect 188822 469338 228266 469574
rect 228502 469338 228586 469574
rect 228822 469338 268266 469574
rect 268502 469338 268586 469574
rect 268822 469338 308266 469574
rect 308502 469338 308586 469574
rect 308822 469338 348266 469574
rect 348502 469338 348586 469574
rect 348822 469338 388266 469574
rect 388502 469338 388586 469574
rect 388822 469338 428266 469574
rect 428502 469338 428586 469574
rect 428822 469338 468266 469574
rect 468502 469338 468586 469574
rect 468822 469338 508266 469574
rect 508502 469338 508586 469574
rect 508822 469338 548266 469574
rect 548502 469338 548586 469574
rect 548822 469338 590142 469574
rect 590378 469338 590462 469574
rect 590698 469338 590730 469574
rect -6806 469306 590730 469338
rect -4886 466174 588810 466206
rect -4886 465938 -4854 466174
rect -4618 465938 -4534 466174
rect -4298 465938 24546 466174
rect 24782 465938 24866 466174
rect 25102 465938 64546 466174
rect 64782 465938 64866 466174
rect 65102 465938 104546 466174
rect 104782 465938 104866 466174
rect 105102 465938 144546 466174
rect 144782 465938 144866 466174
rect 145102 465938 184546 466174
rect 184782 465938 184866 466174
rect 185102 465938 224546 466174
rect 224782 465938 224866 466174
rect 225102 465938 264546 466174
rect 264782 465938 264866 466174
rect 265102 465938 304546 466174
rect 304782 465938 304866 466174
rect 305102 465938 344546 466174
rect 344782 465938 344866 466174
rect 345102 465938 384546 466174
rect 384782 465938 384866 466174
rect 385102 465938 424546 466174
rect 424782 465938 424866 466174
rect 425102 465938 464546 466174
rect 464782 465938 464866 466174
rect 465102 465938 504546 466174
rect 504782 465938 504866 466174
rect 505102 465938 544546 466174
rect 544782 465938 544866 466174
rect 545102 465938 588222 466174
rect 588458 465938 588542 466174
rect 588778 465938 588810 466174
rect -4886 465854 588810 465938
rect -4886 465618 -4854 465854
rect -4618 465618 -4534 465854
rect -4298 465618 24546 465854
rect 24782 465618 24866 465854
rect 25102 465618 64546 465854
rect 64782 465618 64866 465854
rect 65102 465618 104546 465854
rect 104782 465618 104866 465854
rect 105102 465618 144546 465854
rect 144782 465618 144866 465854
rect 145102 465618 184546 465854
rect 184782 465618 184866 465854
rect 185102 465618 224546 465854
rect 224782 465618 224866 465854
rect 225102 465618 264546 465854
rect 264782 465618 264866 465854
rect 265102 465618 304546 465854
rect 304782 465618 304866 465854
rect 305102 465618 344546 465854
rect 344782 465618 344866 465854
rect 345102 465618 384546 465854
rect 384782 465618 384866 465854
rect 385102 465618 424546 465854
rect 424782 465618 424866 465854
rect 425102 465618 464546 465854
rect 464782 465618 464866 465854
rect 465102 465618 504546 465854
rect 504782 465618 504866 465854
rect 505102 465618 544546 465854
rect 544782 465618 544866 465854
rect 545102 465618 588222 465854
rect 588458 465618 588542 465854
rect 588778 465618 588810 465854
rect -4886 465586 588810 465618
rect -2966 462454 586890 462486
rect -2966 462218 -2934 462454
rect -2698 462218 -2614 462454
rect -2378 462218 20826 462454
rect 21062 462218 21146 462454
rect 21382 462218 60826 462454
rect 61062 462218 61146 462454
rect 61382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 140826 462454
rect 141062 462218 141146 462454
rect 141382 462218 180826 462454
rect 181062 462218 181146 462454
rect 181382 462218 220826 462454
rect 221062 462218 221146 462454
rect 221382 462218 260826 462454
rect 261062 462218 261146 462454
rect 261382 462218 300826 462454
rect 301062 462218 301146 462454
rect 301382 462218 340826 462454
rect 341062 462218 341146 462454
rect 341382 462218 380826 462454
rect 381062 462218 381146 462454
rect 381382 462218 420826 462454
rect 421062 462218 421146 462454
rect 421382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 500826 462454
rect 501062 462218 501146 462454
rect 501382 462218 540826 462454
rect 541062 462218 541146 462454
rect 541382 462218 580826 462454
rect 581062 462218 581146 462454
rect 581382 462218 586302 462454
rect 586538 462218 586622 462454
rect 586858 462218 586890 462454
rect -2966 462134 586890 462218
rect -2966 461898 -2934 462134
rect -2698 461898 -2614 462134
rect -2378 461898 20826 462134
rect 21062 461898 21146 462134
rect 21382 461898 60826 462134
rect 61062 461898 61146 462134
rect 61382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 140826 462134
rect 141062 461898 141146 462134
rect 141382 461898 180826 462134
rect 181062 461898 181146 462134
rect 181382 461898 220826 462134
rect 221062 461898 221146 462134
rect 221382 461898 260826 462134
rect 261062 461898 261146 462134
rect 261382 461898 300826 462134
rect 301062 461898 301146 462134
rect 301382 461898 340826 462134
rect 341062 461898 341146 462134
rect 341382 461898 380826 462134
rect 381062 461898 381146 462134
rect 381382 461898 420826 462134
rect 421062 461898 421146 462134
rect 421382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 500826 462134
rect 501062 461898 501146 462134
rect 501382 461898 540826 462134
rect 541062 461898 541146 462134
rect 541382 461898 580826 462134
rect 581062 461898 581146 462134
rect 581382 461898 586302 462134
rect 586538 461898 586622 462134
rect 586858 461898 586890 462134
rect -2966 461866 586890 461898
rect -8726 453614 592650 453646
rect -8726 453378 -7734 453614
rect -7498 453378 -7414 453614
rect -7178 453378 11986 453614
rect 12222 453378 12306 453614
rect 12542 453378 51986 453614
rect 52222 453378 52306 453614
rect 52542 453378 91986 453614
rect 92222 453378 92306 453614
rect 92542 453378 131986 453614
rect 132222 453378 132306 453614
rect 132542 453378 171986 453614
rect 172222 453378 172306 453614
rect 172542 453378 211986 453614
rect 212222 453378 212306 453614
rect 212542 453378 251986 453614
rect 252222 453378 252306 453614
rect 252542 453378 291986 453614
rect 292222 453378 292306 453614
rect 292542 453378 331986 453614
rect 332222 453378 332306 453614
rect 332542 453378 371986 453614
rect 372222 453378 372306 453614
rect 372542 453378 411986 453614
rect 412222 453378 412306 453614
rect 412542 453378 451986 453614
rect 452222 453378 452306 453614
rect 452542 453378 491986 453614
rect 492222 453378 492306 453614
rect 492542 453378 531986 453614
rect 532222 453378 532306 453614
rect 532542 453378 571986 453614
rect 572222 453378 572306 453614
rect 572542 453378 591102 453614
rect 591338 453378 591422 453614
rect 591658 453378 592650 453614
rect -8726 453294 592650 453378
rect -8726 453058 -7734 453294
rect -7498 453058 -7414 453294
rect -7178 453058 11986 453294
rect 12222 453058 12306 453294
rect 12542 453058 51986 453294
rect 52222 453058 52306 453294
rect 52542 453058 91986 453294
rect 92222 453058 92306 453294
rect 92542 453058 131986 453294
rect 132222 453058 132306 453294
rect 132542 453058 171986 453294
rect 172222 453058 172306 453294
rect 172542 453058 211986 453294
rect 212222 453058 212306 453294
rect 212542 453058 251986 453294
rect 252222 453058 252306 453294
rect 252542 453058 291986 453294
rect 292222 453058 292306 453294
rect 292542 453058 331986 453294
rect 332222 453058 332306 453294
rect 332542 453058 371986 453294
rect 372222 453058 372306 453294
rect 372542 453058 411986 453294
rect 412222 453058 412306 453294
rect 412542 453058 451986 453294
rect 452222 453058 452306 453294
rect 452542 453058 491986 453294
rect 492222 453058 492306 453294
rect 492542 453058 531986 453294
rect 532222 453058 532306 453294
rect 532542 453058 571986 453294
rect 572222 453058 572306 453294
rect 572542 453058 591102 453294
rect 591338 453058 591422 453294
rect 591658 453058 592650 453294
rect -8726 453026 592650 453058
rect -6806 449894 590730 449926
rect -6806 449658 -5814 449894
rect -5578 449658 -5494 449894
rect -5258 449658 8266 449894
rect 8502 449658 8586 449894
rect 8822 449658 48266 449894
rect 48502 449658 48586 449894
rect 48822 449658 88266 449894
rect 88502 449658 88586 449894
rect 88822 449658 128266 449894
rect 128502 449658 128586 449894
rect 128822 449658 168266 449894
rect 168502 449658 168586 449894
rect 168822 449658 208266 449894
rect 208502 449658 208586 449894
rect 208822 449658 248266 449894
rect 248502 449658 248586 449894
rect 248822 449658 288266 449894
rect 288502 449658 288586 449894
rect 288822 449658 328266 449894
rect 328502 449658 328586 449894
rect 328822 449658 368266 449894
rect 368502 449658 368586 449894
rect 368822 449658 408266 449894
rect 408502 449658 408586 449894
rect 408822 449658 448266 449894
rect 448502 449658 448586 449894
rect 448822 449658 488266 449894
rect 488502 449658 488586 449894
rect 488822 449658 528266 449894
rect 528502 449658 528586 449894
rect 528822 449658 568266 449894
rect 568502 449658 568586 449894
rect 568822 449658 589182 449894
rect 589418 449658 589502 449894
rect 589738 449658 590730 449894
rect -6806 449574 590730 449658
rect -6806 449338 -5814 449574
rect -5578 449338 -5494 449574
rect -5258 449338 8266 449574
rect 8502 449338 8586 449574
rect 8822 449338 48266 449574
rect 48502 449338 48586 449574
rect 48822 449338 88266 449574
rect 88502 449338 88586 449574
rect 88822 449338 128266 449574
rect 128502 449338 128586 449574
rect 128822 449338 168266 449574
rect 168502 449338 168586 449574
rect 168822 449338 208266 449574
rect 208502 449338 208586 449574
rect 208822 449338 248266 449574
rect 248502 449338 248586 449574
rect 248822 449338 288266 449574
rect 288502 449338 288586 449574
rect 288822 449338 328266 449574
rect 328502 449338 328586 449574
rect 328822 449338 368266 449574
rect 368502 449338 368586 449574
rect 368822 449338 408266 449574
rect 408502 449338 408586 449574
rect 408822 449338 448266 449574
rect 448502 449338 448586 449574
rect 448822 449338 488266 449574
rect 488502 449338 488586 449574
rect 488822 449338 528266 449574
rect 528502 449338 528586 449574
rect 528822 449338 568266 449574
rect 568502 449338 568586 449574
rect 568822 449338 589182 449574
rect 589418 449338 589502 449574
rect 589738 449338 590730 449574
rect -6806 449306 590730 449338
rect -4886 446174 588810 446206
rect -4886 445938 -3894 446174
rect -3658 445938 -3574 446174
rect -3338 445938 4546 446174
rect 4782 445938 4866 446174
rect 5102 445938 44546 446174
rect 44782 445938 44866 446174
rect 45102 445938 84546 446174
rect 84782 445938 84866 446174
rect 85102 445938 124546 446174
rect 124782 445938 124866 446174
rect 125102 445938 164546 446174
rect 164782 445938 164866 446174
rect 165102 445938 204546 446174
rect 204782 445938 204866 446174
rect 205102 445938 244546 446174
rect 244782 445938 244866 446174
rect 245102 445938 284546 446174
rect 284782 445938 284866 446174
rect 285102 445938 324546 446174
rect 324782 445938 324866 446174
rect 325102 445938 364546 446174
rect 364782 445938 364866 446174
rect 365102 445938 404546 446174
rect 404782 445938 404866 446174
rect 405102 445938 444546 446174
rect 444782 445938 444866 446174
rect 445102 445938 484546 446174
rect 484782 445938 484866 446174
rect 485102 445938 524546 446174
rect 524782 445938 524866 446174
rect 525102 445938 564546 446174
rect 564782 445938 564866 446174
rect 565102 445938 587262 446174
rect 587498 445938 587582 446174
rect 587818 445938 588810 446174
rect -4886 445854 588810 445938
rect -4886 445618 -3894 445854
rect -3658 445618 -3574 445854
rect -3338 445618 4546 445854
rect 4782 445618 4866 445854
rect 5102 445618 44546 445854
rect 44782 445618 44866 445854
rect 45102 445618 84546 445854
rect 84782 445618 84866 445854
rect 85102 445618 124546 445854
rect 124782 445618 124866 445854
rect 125102 445618 164546 445854
rect 164782 445618 164866 445854
rect 165102 445618 204546 445854
rect 204782 445618 204866 445854
rect 205102 445618 244546 445854
rect 244782 445618 244866 445854
rect 245102 445618 284546 445854
rect 284782 445618 284866 445854
rect 285102 445618 324546 445854
rect 324782 445618 324866 445854
rect 325102 445618 364546 445854
rect 364782 445618 364866 445854
rect 365102 445618 404546 445854
rect 404782 445618 404866 445854
rect 405102 445618 444546 445854
rect 444782 445618 444866 445854
rect 445102 445618 484546 445854
rect 484782 445618 484866 445854
rect 485102 445618 524546 445854
rect 524782 445618 524866 445854
rect 525102 445618 564546 445854
rect 564782 445618 564866 445854
rect 565102 445618 587262 445854
rect 587498 445618 587582 445854
rect 587818 445618 588810 445854
rect -4886 445586 588810 445618
rect -2966 442454 586890 442486
rect -2966 442218 -1974 442454
rect -1738 442218 -1654 442454
rect -1418 442218 826 442454
rect 1062 442218 1146 442454
rect 1382 442218 40826 442454
rect 41062 442218 41146 442454
rect 41382 442218 80826 442454
rect 81062 442218 81146 442454
rect 81382 442218 120826 442454
rect 121062 442218 121146 442454
rect 121382 442218 160826 442454
rect 161062 442218 161146 442454
rect 161382 442218 200826 442454
rect 201062 442218 201146 442454
rect 201382 442218 240826 442454
rect 241062 442218 241146 442454
rect 241382 442218 280826 442454
rect 281062 442218 281146 442454
rect 281382 442218 320826 442454
rect 321062 442218 321146 442454
rect 321382 442218 360826 442454
rect 361062 442218 361146 442454
rect 361382 442218 400826 442454
rect 401062 442218 401146 442454
rect 401382 442218 440826 442454
rect 441062 442218 441146 442454
rect 441382 442218 480826 442454
rect 481062 442218 481146 442454
rect 481382 442218 520826 442454
rect 521062 442218 521146 442454
rect 521382 442218 560826 442454
rect 561062 442218 561146 442454
rect 561382 442218 585342 442454
rect 585578 442218 585662 442454
rect 585898 442218 586890 442454
rect -2966 442134 586890 442218
rect -2966 441898 -1974 442134
rect -1738 441898 -1654 442134
rect -1418 441898 826 442134
rect 1062 441898 1146 442134
rect 1382 441898 40826 442134
rect 41062 441898 41146 442134
rect 41382 441898 80826 442134
rect 81062 441898 81146 442134
rect 81382 441898 120826 442134
rect 121062 441898 121146 442134
rect 121382 441898 160826 442134
rect 161062 441898 161146 442134
rect 161382 441898 200826 442134
rect 201062 441898 201146 442134
rect 201382 441898 240826 442134
rect 241062 441898 241146 442134
rect 241382 441898 280826 442134
rect 281062 441898 281146 442134
rect 281382 441898 320826 442134
rect 321062 441898 321146 442134
rect 321382 441898 360826 442134
rect 361062 441898 361146 442134
rect 361382 441898 400826 442134
rect 401062 441898 401146 442134
rect 401382 441898 440826 442134
rect 441062 441898 441146 442134
rect 441382 441898 480826 442134
rect 481062 441898 481146 442134
rect 481382 441898 520826 442134
rect 521062 441898 521146 442134
rect 521382 441898 560826 442134
rect 561062 441898 561146 442134
rect 561382 441898 585342 442134
rect 585578 441898 585662 442134
rect 585898 441898 586890 442134
rect -2966 441866 586890 441898
rect -8726 433614 592650 433646
rect -8726 433378 -8694 433614
rect -8458 433378 -8374 433614
rect -8138 433378 31986 433614
rect 32222 433378 32306 433614
rect 32542 433378 71986 433614
rect 72222 433378 72306 433614
rect 72542 433378 111986 433614
rect 112222 433378 112306 433614
rect 112542 433378 151986 433614
rect 152222 433378 152306 433614
rect 152542 433378 191986 433614
rect 192222 433378 192306 433614
rect 192542 433378 231986 433614
rect 232222 433378 232306 433614
rect 232542 433378 271986 433614
rect 272222 433378 272306 433614
rect 272542 433378 311986 433614
rect 312222 433378 312306 433614
rect 312542 433378 351986 433614
rect 352222 433378 352306 433614
rect 352542 433378 391986 433614
rect 392222 433378 392306 433614
rect 392542 433378 431986 433614
rect 432222 433378 432306 433614
rect 432542 433378 471986 433614
rect 472222 433378 472306 433614
rect 472542 433378 511986 433614
rect 512222 433378 512306 433614
rect 512542 433378 551986 433614
rect 552222 433378 552306 433614
rect 552542 433378 592062 433614
rect 592298 433378 592382 433614
rect 592618 433378 592650 433614
rect -8726 433294 592650 433378
rect -8726 433058 -8694 433294
rect -8458 433058 -8374 433294
rect -8138 433058 31986 433294
rect 32222 433058 32306 433294
rect 32542 433058 71986 433294
rect 72222 433058 72306 433294
rect 72542 433058 111986 433294
rect 112222 433058 112306 433294
rect 112542 433058 151986 433294
rect 152222 433058 152306 433294
rect 152542 433058 191986 433294
rect 192222 433058 192306 433294
rect 192542 433058 231986 433294
rect 232222 433058 232306 433294
rect 232542 433058 271986 433294
rect 272222 433058 272306 433294
rect 272542 433058 311986 433294
rect 312222 433058 312306 433294
rect 312542 433058 351986 433294
rect 352222 433058 352306 433294
rect 352542 433058 391986 433294
rect 392222 433058 392306 433294
rect 392542 433058 431986 433294
rect 432222 433058 432306 433294
rect 432542 433058 471986 433294
rect 472222 433058 472306 433294
rect 472542 433058 511986 433294
rect 512222 433058 512306 433294
rect 512542 433058 551986 433294
rect 552222 433058 552306 433294
rect 552542 433058 592062 433294
rect 592298 433058 592382 433294
rect 592618 433058 592650 433294
rect -8726 433026 592650 433058
rect -6806 429894 590730 429926
rect -6806 429658 -6774 429894
rect -6538 429658 -6454 429894
rect -6218 429658 28266 429894
rect 28502 429658 28586 429894
rect 28822 429658 68266 429894
rect 68502 429658 68586 429894
rect 68822 429658 108266 429894
rect 108502 429658 108586 429894
rect 108822 429658 148266 429894
rect 148502 429658 148586 429894
rect 148822 429658 188266 429894
rect 188502 429658 188586 429894
rect 188822 429658 228266 429894
rect 228502 429658 228586 429894
rect 228822 429658 268266 429894
rect 268502 429658 268586 429894
rect 268822 429658 308266 429894
rect 308502 429658 308586 429894
rect 308822 429658 348266 429894
rect 348502 429658 348586 429894
rect 348822 429658 388266 429894
rect 388502 429658 388586 429894
rect 388822 429658 428266 429894
rect 428502 429658 428586 429894
rect 428822 429658 468266 429894
rect 468502 429658 468586 429894
rect 468822 429658 508266 429894
rect 508502 429658 508586 429894
rect 508822 429658 548266 429894
rect 548502 429658 548586 429894
rect 548822 429658 590142 429894
rect 590378 429658 590462 429894
rect 590698 429658 590730 429894
rect -6806 429574 590730 429658
rect -6806 429338 -6774 429574
rect -6538 429338 -6454 429574
rect -6218 429338 28266 429574
rect 28502 429338 28586 429574
rect 28822 429338 68266 429574
rect 68502 429338 68586 429574
rect 68822 429338 108266 429574
rect 108502 429338 108586 429574
rect 108822 429338 148266 429574
rect 148502 429338 148586 429574
rect 148822 429338 188266 429574
rect 188502 429338 188586 429574
rect 188822 429338 228266 429574
rect 228502 429338 228586 429574
rect 228822 429338 268266 429574
rect 268502 429338 268586 429574
rect 268822 429338 308266 429574
rect 308502 429338 308586 429574
rect 308822 429338 348266 429574
rect 348502 429338 348586 429574
rect 348822 429338 388266 429574
rect 388502 429338 388586 429574
rect 388822 429338 428266 429574
rect 428502 429338 428586 429574
rect 428822 429338 468266 429574
rect 468502 429338 468586 429574
rect 468822 429338 508266 429574
rect 508502 429338 508586 429574
rect 508822 429338 548266 429574
rect 548502 429338 548586 429574
rect 548822 429338 590142 429574
rect 590378 429338 590462 429574
rect 590698 429338 590730 429574
rect -6806 429306 590730 429338
rect -4886 426174 588810 426206
rect -4886 425938 -4854 426174
rect -4618 425938 -4534 426174
rect -4298 425938 24546 426174
rect 24782 425938 24866 426174
rect 25102 425938 64546 426174
rect 64782 425938 64866 426174
rect 65102 425938 104546 426174
rect 104782 425938 104866 426174
rect 105102 425938 144546 426174
rect 144782 425938 144866 426174
rect 145102 425938 184546 426174
rect 184782 425938 184866 426174
rect 185102 425938 224546 426174
rect 224782 425938 224866 426174
rect 225102 425938 264546 426174
rect 264782 425938 264866 426174
rect 265102 425938 304546 426174
rect 304782 425938 304866 426174
rect 305102 425938 344546 426174
rect 344782 425938 344866 426174
rect 345102 425938 384546 426174
rect 384782 425938 384866 426174
rect 385102 425938 424546 426174
rect 424782 425938 424866 426174
rect 425102 425938 464546 426174
rect 464782 425938 464866 426174
rect 465102 425938 504546 426174
rect 504782 425938 504866 426174
rect 505102 425938 544546 426174
rect 544782 425938 544866 426174
rect 545102 425938 588222 426174
rect 588458 425938 588542 426174
rect 588778 425938 588810 426174
rect -4886 425854 588810 425938
rect -4886 425618 -4854 425854
rect -4618 425618 -4534 425854
rect -4298 425618 24546 425854
rect 24782 425618 24866 425854
rect 25102 425618 64546 425854
rect 64782 425618 64866 425854
rect 65102 425618 104546 425854
rect 104782 425618 104866 425854
rect 105102 425618 144546 425854
rect 144782 425618 144866 425854
rect 145102 425618 184546 425854
rect 184782 425618 184866 425854
rect 185102 425618 224546 425854
rect 224782 425618 224866 425854
rect 225102 425618 264546 425854
rect 264782 425618 264866 425854
rect 265102 425618 304546 425854
rect 304782 425618 304866 425854
rect 305102 425618 344546 425854
rect 344782 425618 344866 425854
rect 345102 425618 384546 425854
rect 384782 425618 384866 425854
rect 385102 425618 424546 425854
rect 424782 425618 424866 425854
rect 425102 425618 464546 425854
rect 464782 425618 464866 425854
rect 465102 425618 504546 425854
rect 504782 425618 504866 425854
rect 505102 425618 544546 425854
rect 544782 425618 544866 425854
rect 545102 425618 588222 425854
rect 588458 425618 588542 425854
rect 588778 425618 588810 425854
rect -4886 425586 588810 425618
rect -2966 422454 586890 422486
rect -2966 422218 -2934 422454
rect -2698 422218 -2614 422454
rect -2378 422218 20826 422454
rect 21062 422218 21146 422454
rect 21382 422218 60826 422454
rect 61062 422218 61146 422454
rect 61382 422218 100826 422454
rect 101062 422218 101146 422454
rect 101382 422218 140826 422454
rect 141062 422218 141146 422454
rect 141382 422218 180826 422454
rect 181062 422218 181146 422454
rect 181382 422218 220826 422454
rect 221062 422218 221146 422454
rect 221382 422218 260826 422454
rect 261062 422218 261146 422454
rect 261382 422218 300826 422454
rect 301062 422218 301146 422454
rect 301382 422218 340826 422454
rect 341062 422218 341146 422454
rect 341382 422218 380826 422454
rect 381062 422218 381146 422454
rect 381382 422218 420826 422454
rect 421062 422218 421146 422454
rect 421382 422218 460826 422454
rect 461062 422218 461146 422454
rect 461382 422218 500826 422454
rect 501062 422218 501146 422454
rect 501382 422218 540826 422454
rect 541062 422218 541146 422454
rect 541382 422218 580826 422454
rect 581062 422218 581146 422454
rect 581382 422218 586302 422454
rect 586538 422218 586622 422454
rect 586858 422218 586890 422454
rect -2966 422134 586890 422218
rect -2966 421898 -2934 422134
rect -2698 421898 -2614 422134
rect -2378 421898 20826 422134
rect 21062 421898 21146 422134
rect 21382 421898 60826 422134
rect 61062 421898 61146 422134
rect 61382 421898 100826 422134
rect 101062 421898 101146 422134
rect 101382 421898 140826 422134
rect 141062 421898 141146 422134
rect 141382 421898 180826 422134
rect 181062 421898 181146 422134
rect 181382 421898 220826 422134
rect 221062 421898 221146 422134
rect 221382 421898 260826 422134
rect 261062 421898 261146 422134
rect 261382 421898 300826 422134
rect 301062 421898 301146 422134
rect 301382 421898 340826 422134
rect 341062 421898 341146 422134
rect 341382 421898 380826 422134
rect 381062 421898 381146 422134
rect 381382 421898 420826 422134
rect 421062 421898 421146 422134
rect 421382 421898 460826 422134
rect 461062 421898 461146 422134
rect 461382 421898 500826 422134
rect 501062 421898 501146 422134
rect 501382 421898 540826 422134
rect 541062 421898 541146 422134
rect 541382 421898 580826 422134
rect 581062 421898 581146 422134
rect 581382 421898 586302 422134
rect 586538 421898 586622 422134
rect 586858 421898 586890 422134
rect -2966 421866 586890 421898
rect -8726 413614 592650 413646
rect -8726 413378 -7734 413614
rect -7498 413378 -7414 413614
rect -7178 413378 11986 413614
rect 12222 413378 12306 413614
rect 12542 413378 51986 413614
rect 52222 413378 52306 413614
rect 52542 413378 91986 413614
rect 92222 413378 92306 413614
rect 92542 413378 131986 413614
rect 132222 413378 132306 413614
rect 132542 413378 171986 413614
rect 172222 413378 172306 413614
rect 172542 413378 211986 413614
rect 212222 413378 212306 413614
rect 212542 413378 251986 413614
rect 252222 413378 252306 413614
rect 252542 413378 291986 413614
rect 292222 413378 292306 413614
rect 292542 413378 331986 413614
rect 332222 413378 332306 413614
rect 332542 413378 371986 413614
rect 372222 413378 372306 413614
rect 372542 413378 411986 413614
rect 412222 413378 412306 413614
rect 412542 413378 451986 413614
rect 452222 413378 452306 413614
rect 452542 413378 491986 413614
rect 492222 413378 492306 413614
rect 492542 413378 531986 413614
rect 532222 413378 532306 413614
rect 532542 413378 571986 413614
rect 572222 413378 572306 413614
rect 572542 413378 591102 413614
rect 591338 413378 591422 413614
rect 591658 413378 592650 413614
rect -8726 413294 592650 413378
rect -8726 413058 -7734 413294
rect -7498 413058 -7414 413294
rect -7178 413058 11986 413294
rect 12222 413058 12306 413294
rect 12542 413058 51986 413294
rect 52222 413058 52306 413294
rect 52542 413058 91986 413294
rect 92222 413058 92306 413294
rect 92542 413058 131986 413294
rect 132222 413058 132306 413294
rect 132542 413058 171986 413294
rect 172222 413058 172306 413294
rect 172542 413058 211986 413294
rect 212222 413058 212306 413294
rect 212542 413058 251986 413294
rect 252222 413058 252306 413294
rect 252542 413058 291986 413294
rect 292222 413058 292306 413294
rect 292542 413058 331986 413294
rect 332222 413058 332306 413294
rect 332542 413058 371986 413294
rect 372222 413058 372306 413294
rect 372542 413058 411986 413294
rect 412222 413058 412306 413294
rect 412542 413058 451986 413294
rect 452222 413058 452306 413294
rect 452542 413058 491986 413294
rect 492222 413058 492306 413294
rect 492542 413058 531986 413294
rect 532222 413058 532306 413294
rect 532542 413058 571986 413294
rect 572222 413058 572306 413294
rect 572542 413058 591102 413294
rect 591338 413058 591422 413294
rect 591658 413058 592650 413294
rect -8726 413026 592650 413058
rect -6806 409894 590730 409926
rect -6806 409658 -5814 409894
rect -5578 409658 -5494 409894
rect -5258 409658 8266 409894
rect 8502 409658 8586 409894
rect 8822 409658 48266 409894
rect 48502 409658 48586 409894
rect 48822 409658 88266 409894
rect 88502 409658 88586 409894
rect 88822 409658 128266 409894
rect 128502 409658 128586 409894
rect 128822 409658 168266 409894
rect 168502 409658 168586 409894
rect 168822 409658 208266 409894
rect 208502 409658 208586 409894
rect 208822 409658 248266 409894
rect 248502 409658 248586 409894
rect 248822 409658 288266 409894
rect 288502 409658 288586 409894
rect 288822 409658 328266 409894
rect 328502 409658 328586 409894
rect 328822 409658 368266 409894
rect 368502 409658 368586 409894
rect 368822 409658 408266 409894
rect 408502 409658 408586 409894
rect 408822 409658 448266 409894
rect 448502 409658 448586 409894
rect 448822 409658 488266 409894
rect 488502 409658 488586 409894
rect 488822 409658 528266 409894
rect 528502 409658 528586 409894
rect 528822 409658 568266 409894
rect 568502 409658 568586 409894
rect 568822 409658 589182 409894
rect 589418 409658 589502 409894
rect 589738 409658 590730 409894
rect -6806 409574 590730 409658
rect -6806 409338 -5814 409574
rect -5578 409338 -5494 409574
rect -5258 409338 8266 409574
rect 8502 409338 8586 409574
rect 8822 409338 48266 409574
rect 48502 409338 48586 409574
rect 48822 409338 88266 409574
rect 88502 409338 88586 409574
rect 88822 409338 128266 409574
rect 128502 409338 128586 409574
rect 128822 409338 168266 409574
rect 168502 409338 168586 409574
rect 168822 409338 208266 409574
rect 208502 409338 208586 409574
rect 208822 409338 248266 409574
rect 248502 409338 248586 409574
rect 248822 409338 288266 409574
rect 288502 409338 288586 409574
rect 288822 409338 328266 409574
rect 328502 409338 328586 409574
rect 328822 409338 368266 409574
rect 368502 409338 368586 409574
rect 368822 409338 408266 409574
rect 408502 409338 408586 409574
rect 408822 409338 448266 409574
rect 448502 409338 448586 409574
rect 448822 409338 488266 409574
rect 488502 409338 488586 409574
rect 488822 409338 528266 409574
rect 528502 409338 528586 409574
rect 528822 409338 568266 409574
rect 568502 409338 568586 409574
rect 568822 409338 589182 409574
rect 589418 409338 589502 409574
rect 589738 409338 590730 409574
rect -6806 409306 590730 409338
rect -4886 406174 588810 406206
rect -4886 405938 -3894 406174
rect -3658 405938 -3574 406174
rect -3338 405938 4546 406174
rect 4782 405938 4866 406174
rect 5102 405938 44546 406174
rect 44782 405938 44866 406174
rect 45102 405938 84546 406174
rect 84782 405938 84866 406174
rect 85102 405938 124546 406174
rect 124782 405938 124866 406174
rect 125102 405938 164546 406174
rect 164782 405938 164866 406174
rect 165102 405938 204546 406174
rect 204782 405938 204866 406174
rect 205102 405938 244546 406174
rect 244782 405938 244866 406174
rect 245102 405938 284546 406174
rect 284782 405938 284866 406174
rect 285102 405938 324546 406174
rect 324782 405938 324866 406174
rect 325102 405938 364546 406174
rect 364782 405938 364866 406174
rect 365102 405938 404546 406174
rect 404782 405938 404866 406174
rect 405102 405938 444546 406174
rect 444782 405938 444866 406174
rect 445102 405938 484546 406174
rect 484782 405938 484866 406174
rect 485102 405938 524546 406174
rect 524782 405938 524866 406174
rect 525102 405938 564546 406174
rect 564782 405938 564866 406174
rect 565102 405938 587262 406174
rect 587498 405938 587582 406174
rect 587818 405938 588810 406174
rect -4886 405854 588810 405938
rect -4886 405618 -3894 405854
rect -3658 405618 -3574 405854
rect -3338 405618 4546 405854
rect 4782 405618 4866 405854
rect 5102 405618 44546 405854
rect 44782 405618 44866 405854
rect 45102 405618 84546 405854
rect 84782 405618 84866 405854
rect 85102 405618 124546 405854
rect 124782 405618 124866 405854
rect 125102 405618 164546 405854
rect 164782 405618 164866 405854
rect 165102 405618 204546 405854
rect 204782 405618 204866 405854
rect 205102 405618 244546 405854
rect 244782 405618 244866 405854
rect 245102 405618 284546 405854
rect 284782 405618 284866 405854
rect 285102 405618 324546 405854
rect 324782 405618 324866 405854
rect 325102 405618 364546 405854
rect 364782 405618 364866 405854
rect 365102 405618 404546 405854
rect 404782 405618 404866 405854
rect 405102 405618 444546 405854
rect 444782 405618 444866 405854
rect 445102 405618 484546 405854
rect 484782 405618 484866 405854
rect 485102 405618 524546 405854
rect 524782 405618 524866 405854
rect 525102 405618 564546 405854
rect 564782 405618 564866 405854
rect 565102 405618 587262 405854
rect 587498 405618 587582 405854
rect 587818 405618 588810 405854
rect -4886 405586 588810 405618
rect -2966 402454 586890 402486
rect -2966 402218 -1974 402454
rect -1738 402218 -1654 402454
rect -1418 402218 826 402454
rect 1062 402218 1146 402454
rect 1382 402218 40826 402454
rect 41062 402218 41146 402454
rect 41382 402218 80826 402454
rect 81062 402218 81146 402454
rect 81382 402218 120826 402454
rect 121062 402218 121146 402454
rect 121382 402218 160826 402454
rect 161062 402218 161146 402454
rect 161382 402218 200826 402454
rect 201062 402218 201146 402454
rect 201382 402218 240826 402454
rect 241062 402218 241146 402454
rect 241382 402218 280826 402454
rect 281062 402218 281146 402454
rect 281382 402218 320826 402454
rect 321062 402218 321146 402454
rect 321382 402218 360826 402454
rect 361062 402218 361146 402454
rect 361382 402218 400826 402454
rect 401062 402218 401146 402454
rect 401382 402218 440826 402454
rect 441062 402218 441146 402454
rect 441382 402218 480826 402454
rect 481062 402218 481146 402454
rect 481382 402218 520826 402454
rect 521062 402218 521146 402454
rect 521382 402218 560826 402454
rect 561062 402218 561146 402454
rect 561382 402218 585342 402454
rect 585578 402218 585662 402454
rect 585898 402218 586890 402454
rect -2966 402134 586890 402218
rect -2966 401898 -1974 402134
rect -1738 401898 -1654 402134
rect -1418 401898 826 402134
rect 1062 401898 1146 402134
rect 1382 401898 40826 402134
rect 41062 401898 41146 402134
rect 41382 401898 80826 402134
rect 81062 401898 81146 402134
rect 81382 401898 120826 402134
rect 121062 401898 121146 402134
rect 121382 401898 160826 402134
rect 161062 401898 161146 402134
rect 161382 401898 200826 402134
rect 201062 401898 201146 402134
rect 201382 401898 240826 402134
rect 241062 401898 241146 402134
rect 241382 401898 280826 402134
rect 281062 401898 281146 402134
rect 281382 401898 320826 402134
rect 321062 401898 321146 402134
rect 321382 401898 360826 402134
rect 361062 401898 361146 402134
rect 361382 401898 400826 402134
rect 401062 401898 401146 402134
rect 401382 401898 440826 402134
rect 441062 401898 441146 402134
rect 441382 401898 480826 402134
rect 481062 401898 481146 402134
rect 481382 401898 520826 402134
rect 521062 401898 521146 402134
rect 521382 401898 560826 402134
rect 561062 401898 561146 402134
rect 561382 401898 585342 402134
rect 585578 401898 585662 402134
rect 585898 401898 586890 402134
rect -2966 401866 586890 401898
rect -8726 393614 592650 393646
rect -8726 393378 -8694 393614
rect -8458 393378 -8374 393614
rect -8138 393378 31986 393614
rect 32222 393378 32306 393614
rect 32542 393378 71986 393614
rect 72222 393378 72306 393614
rect 72542 393378 111986 393614
rect 112222 393378 112306 393614
rect 112542 393378 151986 393614
rect 152222 393378 152306 393614
rect 152542 393378 191986 393614
rect 192222 393378 192306 393614
rect 192542 393378 231986 393614
rect 232222 393378 232306 393614
rect 232542 393378 271986 393614
rect 272222 393378 272306 393614
rect 272542 393378 311986 393614
rect 312222 393378 312306 393614
rect 312542 393378 351986 393614
rect 352222 393378 352306 393614
rect 352542 393378 391986 393614
rect 392222 393378 392306 393614
rect 392542 393378 431986 393614
rect 432222 393378 432306 393614
rect 432542 393378 471986 393614
rect 472222 393378 472306 393614
rect 472542 393378 511986 393614
rect 512222 393378 512306 393614
rect 512542 393378 551986 393614
rect 552222 393378 552306 393614
rect 552542 393378 592062 393614
rect 592298 393378 592382 393614
rect 592618 393378 592650 393614
rect -8726 393294 592650 393378
rect -8726 393058 -8694 393294
rect -8458 393058 -8374 393294
rect -8138 393058 31986 393294
rect 32222 393058 32306 393294
rect 32542 393058 71986 393294
rect 72222 393058 72306 393294
rect 72542 393058 111986 393294
rect 112222 393058 112306 393294
rect 112542 393058 151986 393294
rect 152222 393058 152306 393294
rect 152542 393058 191986 393294
rect 192222 393058 192306 393294
rect 192542 393058 231986 393294
rect 232222 393058 232306 393294
rect 232542 393058 271986 393294
rect 272222 393058 272306 393294
rect 272542 393058 311986 393294
rect 312222 393058 312306 393294
rect 312542 393058 351986 393294
rect 352222 393058 352306 393294
rect 352542 393058 391986 393294
rect 392222 393058 392306 393294
rect 392542 393058 431986 393294
rect 432222 393058 432306 393294
rect 432542 393058 471986 393294
rect 472222 393058 472306 393294
rect 472542 393058 511986 393294
rect 512222 393058 512306 393294
rect 512542 393058 551986 393294
rect 552222 393058 552306 393294
rect 552542 393058 592062 393294
rect 592298 393058 592382 393294
rect 592618 393058 592650 393294
rect -8726 393026 592650 393058
rect -6806 389894 590730 389926
rect -6806 389658 -6774 389894
rect -6538 389658 -6454 389894
rect -6218 389658 28266 389894
rect 28502 389658 28586 389894
rect 28822 389658 68266 389894
rect 68502 389658 68586 389894
rect 68822 389658 108266 389894
rect 108502 389658 108586 389894
rect 108822 389658 148266 389894
rect 148502 389658 148586 389894
rect 148822 389658 188266 389894
rect 188502 389658 188586 389894
rect 188822 389658 228266 389894
rect 228502 389658 228586 389894
rect 228822 389658 268266 389894
rect 268502 389658 268586 389894
rect 268822 389658 308266 389894
rect 308502 389658 308586 389894
rect 308822 389658 348266 389894
rect 348502 389658 348586 389894
rect 348822 389658 388266 389894
rect 388502 389658 388586 389894
rect 388822 389658 428266 389894
rect 428502 389658 428586 389894
rect 428822 389658 468266 389894
rect 468502 389658 468586 389894
rect 468822 389658 508266 389894
rect 508502 389658 508586 389894
rect 508822 389658 548266 389894
rect 548502 389658 548586 389894
rect 548822 389658 590142 389894
rect 590378 389658 590462 389894
rect 590698 389658 590730 389894
rect -6806 389574 590730 389658
rect -6806 389338 -6774 389574
rect -6538 389338 -6454 389574
rect -6218 389338 28266 389574
rect 28502 389338 28586 389574
rect 28822 389338 68266 389574
rect 68502 389338 68586 389574
rect 68822 389338 108266 389574
rect 108502 389338 108586 389574
rect 108822 389338 148266 389574
rect 148502 389338 148586 389574
rect 148822 389338 188266 389574
rect 188502 389338 188586 389574
rect 188822 389338 228266 389574
rect 228502 389338 228586 389574
rect 228822 389338 268266 389574
rect 268502 389338 268586 389574
rect 268822 389338 308266 389574
rect 308502 389338 308586 389574
rect 308822 389338 348266 389574
rect 348502 389338 348586 389574
rect 348822 389338 388266 389574
rect 388502 389338 388586 389574
rect 388822 389338 428266 389574
rect 428502 389338 428586 389574
rect 428822 389338 468266 389574
rect 468502 389338 468586 389574
rect 468822 389338 508266 389574
rect 508502 389338 508586 389574
rect 508822 389338 548266 389574
rect 548502 389338 548586 389574
rect 548822 389338 590142 389574
rect 590378 389338 590462 389574
rect 590698 389338 590730 389574
rect -6806 389306 590730 389338
rect -4886 386174 588810 386206
rect -4886 385938 -4854 386174
rect -4618 385938 -4534 386174
rect -4298 385938 24546 386174
rect 24782 385938 24866 386174
rect 25102 385938 64546 386174
rect 64782 385938 64866 386174
rect 65102 385938 104546 386174
rect 104782 385938 104866 386174
rect 105102 385938 144546 386174
rect 144782 385938 144866 386174
rect 145102 385938 184546 386174
rect 184782 385938 184866 386174
rect 185102 385938 224546 386174
rect 224782 385938 224866 386174
rect 225102 385938 264546 386174
rect 264782 385938 264866 386174
rect 265102 385938 304546 386174
rect 304782 385938 304866 386174
rect 305102 385938 344546 386174
rect 344782 385938 344866 386174
rect 345102 385938 384546 386174
rect 384782 385938 384866 386174
rect 385102 385938 424546 386174
rect 424782 385938 424866 386174
rect 425102 385938 464546 386174
rect 464782 385938 464866 386174
rect 465102 385938 504546 386174
rect 504782 385938 504866 386174
rect 505102 385938 544546 386174
rect 544782 385938 544866 386174
rect 545102 385938 588222 386174
rect 588458 385938 588542 386174
rect 588778 385938 588810 386174
rect -4886 385854 588810 385938
rect -4886 385618 -4854 385854
rect -4618 385618 -4534 385854
rect -4298 385618 24546 385854
rect 24782 385618 24866 385854
rect 25102 385618 64546 385854
rect 64782 385618 64866 385854
rect 65102 385618 104546 385854
rect 104782 385618 104866 385854
rect 105102 385618 144546 385854
rect 144782 385618 144866 385854
rect 145102 385618 184546 385854
rect 184782 385618 184866 385854
rect 185102 385618 224546 385854
rect 224782 385618 224866 385854
rect 225102 385618 264546 385854
rect 264782 385618 264866 385854
rect 265102 385618 304546 385854
rect 304782 385618 304866 385854
rect 305102 385618 344546 385854
rect 344782 385618 344866 385854
rect 345102 385618 384546 385854
rect 384782 385618 384866 385854
rect 385102 385618 424546 385854
rect 424782 385618 424866 385854
rect 425102 385618 464546 385854
rect 464782 385618 464866 385854
rect 465102 385618 504546 385854
rect 504782 385618 504866 385854
rect 505102 385618 544546 385854
rect 544782 385618 544866 385854
rect 545102 385618 588222 385854
rect 588458 385618 588542 385854
rect 588778 385618 588810 385854
rect -4886 385586 588810 385618
rect -2966 382454 586890 382486
rect -2966 382218 -2934 382454
rect -2698 382218 -2614 382454
rect -2378 382218 20826 382454
rect 21062 382218 21146 382454
rect 21382 382218 60826 382454
rect 61062 382218 61146 382454
rect 61382 382218 100826 382454
rect 101062 382218 101146 382454
rect 101382 382218 140826 382454
rect 141062 382218 141146 382454
rect 141382 382218 180826 382454
rect 181062 382218 181146 382454
rect 181382 382218 220826 382454
rect 221062 382218 221146 382454
rect 221382 382218 260826 382454
rect 261062 382218 261146 382454
rect 261382 382218 300826 382454
rect 301062 382218 301146 382454
rect 301382 382218 340826 382454
rect 341062 382218 341146 382454
rect 341382 382218 380826 382454
rect 381062 382218 381146 382454
rect 381382 382218 420826 382454
rect 421062 382218 421146 382454
rect 421382 382218 460826 382454
rect 461062 382218 461146 382454
rect 461382 382218 500826 382454
rect 501062 382218 501146 382454
rect 501382 382218 540826 382454
rect 541062 382218 541146 382454
rect 541382 382218 580826 382454
rect 581062 382218 581146 382454
rect 581382 382218 586302 382454
rect 586538 382218 586622 382454
rect 586858 382218 586890 382454
rect -2966 382134 586890 382218
rect -2966 381898 -2934 382134
rect -2698 381898 -2614 382134
rect -2378 381898 20826 382134
rect 21062 381898 21146 382134
rect 21382 381898 60826 382134
rect 61062 381898 61146 382134
rect 61382 381898 100826 382134
rect 101062 381898 101146 382134
rect 101382 381898 140826 382134
rect 141062 381898 141146 382134
rect 141382 381898 180826 382134
rect 181062 381898 181146 382134
rect 181382 381898 220826 382134
rect 221062 381898 221146 382134
rect 221382 381898 260826 382134
rect 261062 381898 261146 382134
rect 261382 381898 300826 382134
rect 301062 381898 301146 382134
rect 301382 381898 340826 382134
rect 341062 381898 341146 382134
rect 341382 381898 380826 382134
rect 381062 381898 381146 382134
rect 381382 381898 420826 382134
rect 421062 381898 421146 382134
rect 421382 381898 460826 382134
rect 461062 381898 461146 382134
rect 461382 381898 500826 382134
rect 501062 381898 501146 382134
rect 501382 381898 540826 382134
rect 541062 381898 541146 382134
rect 541382 381898 580826 382134
rect 581062 381898 581146 382134
rect 581382 381898 586302 382134
rect 586538 381898 586622 382134
rect 586858 381898 586890 382134
rect -2966 381866 586890 381898
rect -8726 373614 592650 373646
rect -8726 373378 -7734 373614
rect -7498 373378 -7414 373614
rect -7178 373378 11986 373614
rect 12222 373378 12306 373614
rect 12542 373378 51986 373614
rect 52222 373378 52306 373614
rect 52542 373378 91986 373614
rect 92222 373378 92306 373614
rect 92542 373378 131986 373614
rect 132222 373378 132306 373614
rect 132542 373378 171986 373614
rect 172222 373378 172306 373614
rect 172542 373378 211986 373614
rect 212222 373378 212306 373614
rect 212542 373378 251986 373614
rect 252222 373378 252306 373614
rect 252542 373378 291986 373614
rect 292222 373378 292306 373614
rect 292542 373378 331986 373614
rect 332222 373378 332306 373614
rect 332542 373378 371986 373614
rect 372222 373378 372306 373614
rect 372542 373378 411986 373614
rect 412222 373378 412306 373614
rect 412542 373378 451986 373614
rect 452222 373378 452306 373614
rect 452542 373378 491986 373614
rect 492222 373378 492306 373614
rect 492542 373378 531986 373614
rect 532222 373378 532306 373614
rect 532542 373378 571986 373614
rect 572222 373378 572306 373614
rect 572542 373378 591102 373614
rect 591338 373378 591422 373614
rect 591658 373378 592650 373614
rect -8726 373294 592650 373378
rect -8726 373058 -7734 373294
rect -7498 373058 -7414 373294
rect -7178 373058 11986 373294
rect 12222 373058 12306 373294
rect 12542 373058 51986 373294
rect 52222 373058 52306 373294
rect 52542 373058 91986 373294
rect 92222 373058 92306 373294
rect 92542 373058 131986 373294
rect 132222 373058 132306 373294
rect 132542 373058 171986 373294
rect 172222 373058 172306 373294
rect 172542 373058 211986 373294
rect 212222 373058 212306 373294
rect 212542 373058 251986 373294
rect 252222 373058 252306 373294
rect 252542 373058 291986 373294
rect 292222 373058 292306 373294
rect 292542 373058 331986 373294
rect 332222 373058 332306 373294
rect 332542 373058 371986 373294
rect 372222 373058 372306 373294
rect 372542 373058 411986 373294
rect 412222 373058 412306 373294
rect 412542 373058 451986 373294
rect 452222 373058 452306 373294
rect 452542 373058 491986 373294
rect 492222 373058 492306 373294
rect 492542 373058 531986 373294
rect 532222 373058 532306 373294
rect 532542 373058 571986 373294
rect 572222 373058 572306 373294
rect 572542 373058 591102 373294
rect 591338 373058 591422 373294
rect 591658 373058 592650 373294
rect -8726 373026 592650 373058
rect -6806 369894 590730 369926
rect -6806 369658 -5814 369894
rect -5578 369658 -5494 369894
rect -5258 369658 8266 369894
rect 8502 369658 8586 369894
rect 8822 369658 48266 369894
rect 48502 369658 48586 369894
rect 48822 369658 88266 369894
rect 88502 369658 88586 369894
rect 88822 369658 128266 369894
rect 128502 369658 128586 369894
rect 128822 369658 168266 369894
rect 168502 369658 168586 369894
rect 168822 369658 208266 369894
rect 208502 369658 208586 369894
rect 208822 369658 248266 369894
rect 248502 369658 248586 369894
rect 248822 369658 288266 369894
rect 288502 369658 288586 369894
rect 288822 369658 328266 369894
rect 328502 369658 328586 369894
rect 328822 369658 368266 369894
rect 368502 369658 368586 369894
rect 368822 369658 408266 369894
rect 408502 369658 408586 369894
rect 408822 369658 448266 369894
rect 448502 369658 448586 369894
rect 448822 369658 488266 369894
rect 488502 369658 488586 369894
rect 488822 369658 528266 369894
rect 528502 369658 528586 369894
rect 528822 369658 568266 369894
rect 568502 369658 568586 369894
rect 568822 369658 589182 369894
rect 589418 369658 589502 369894
rect 589738 369658 590730 369894
rect -6806 369574 590730 369658
rect -6806 369338 -5814 369574
rect -5578 369338 -5494 369574
rect -5258 369338 8266 369574
rect 8502 369338 8586 369574
rect 8822 369338 48266 369574
rect 48502 369338 48586 369574
rect 48822 369338 88266 369574
rect 88502 369338 88586 369574
rect 88822 369338 128266 369574
rect 128502 369338 128586 369574
rect 128822 369338 168266 369574
rect 168502 369338 168586 369574
rect 168822 369338 208266 369574
rect 208502 369338 208586 369574
rect 208822 369338 248266 369574
rect 248502 369338 248586 369574
rect 248822 369338 288266 369574
rect 288502 369338 288586 369574
rect 288822 369338 328266 369574
rect 328502 369338 328586 369574
rect 328822 369338 368266 369574
rect 368502 369338 368586 369574
rect 368822 369338 408266 369574
rect 408502 369338 408586 369574
rect 408822 369338 448266 369574
rect 448502 369338 448586 369574
rect 448822 369338 488266 369574
rect 488502 369338 488586 369574
rect 488822 369338 528266 369574
rect 528502 369338 528586 369574
rect 528822 369338 568266 369574
rect 568502 369338 568586 369574
rect 568822 369338 589182 369574
rect 589418 369338 589502 369574
rect 589738 369338 590730 369574
rect -6806 369306 590730 369338
rect -4886 366174 588810 366206
rect -4886 365938 -3894 366174
rect -3658 365938 -3574 366174
rect -3338 365938 4546 366174
rect 4782 365938 4866 366174
rect 5102 365938 44546 366174
rect 44782 365938 44866 366174
rect 45102 365938 84546 366174
rect 84782 365938 84866 366174
rect 85102 365938 124546 366174
rect 124782 365938 124866 366174
rect 125102 365938 164546 366174
rect 164782 365938 164866 366174
rect 165102 365938 204546 366174
rect 204782 365938 204866 366174
rect 205102 365938 244546 366174
rect 244782 365938 244866 366174
rect 245102 365938 284546 366174
rect 284782 365938 284866 366174
rect 285102 365938 324546 366174
rect 324782 365938 324866 366174
rect 325102 365938 364546 366174
rect 364782 365938 364866 366174
rect 365102 365938 404546 366174
rect 404782 365938 404866 366174
rect 405102 365938 444546 366174
rect 444782 365938 444866 366174
rect 445102 365938 484546 366174
rect 484782 365938 484866 366174
rect 485102 365938 524546 366174
rect 524782 365938 524866 366174
rect 525102 365938 564546 366174
rect 564782 365938 564866 366174
rect 565102 365938 587262 366174
rect 587498 365938 587582 366174
rect 587818 365938 588810 366174
rect -4886 365854 588810 365938
rect -4886 365618 -3894 365854
rect -3658 365618 -3574 365854
rect -3338 365618 4546 365854
rect 4782 365618 4866 365854
rect 5102 365618 44546 365854
rect 44782 365618 44866 365854
rect 45102 365618 84546 365854
rect 84782 365618 84866 365854
rect 85102 365618 124546 365854
rect 124782 365618 124866 365854
rect 125102 365618 164546 365854
rect 164782 365618 164866 365854
rect 165102 365618 204546 365854
rect 204782 365618 204866 365854
rect 205102 365618 244546 365854
rect 244782 365618 244866 365854
rect 245102 365618 284546 365854
rect 284782 365618 284866 365854
rect 285102 365618 324546 365854
rect 324782 365618 324866 365854
rect 325102 365618 364546 365854
rect 364782 365618 364866 365854
rect 365102 365618 404546 365854
rect 404782 365618 404866 365854
rect 405102 365618 444546 365854
rect 444782 365618 444866 365854
rect 445102 365618 484546 365854
rect 484782 365618 484866 365854
rect 485102 365618 524546 365854
rect 524782 365618 524866 365854
rect 525102 365618 564546 365854
rect 564782 365618 564866 365854
rect 565102 365618 587262 365854
rect 587498 365618 587582 365854
rect 587818 365618 588810 365854
rect -4886 365586 588810 365618
rect -2966 362454 586890 362486
rect -2966 362218 -1974 362454
rect -1738 362218 -1654 362454
rect -1418 362218 826 362454
rect 1062 362218 1146 362454
rect 1382 362218 40826 362454
rect 41062 362218 41146 362454
rect 41382 362218 80826 362454
rect 81062 362218 81146 362454
rect 81382 362218 120826 362454
rect 121062 362218 121146 362454
rect 121382 362218 160826 362454
rect 161062 362218 161146 362454
rect 161382 362218 200826 362454
rect 201062 362218 201146 362454
rect 201382 362218 240826 362454
rect 241062 362218 241146 362454
rect 241382 362218 280826 362454
rect 281062 362218 281146 362454
rect 281382 362218 320826 362454
rect 321062 362218 321146 362454
rect 321382 362218 360826 362454
rect 361062 362218 361146 362454
rect 361382 362218 400826 362454
rect 401062 362218 401146 362454
rect 401382 362218 440826 362454
rect 441062 362218 441146 362454
rect 441382 362218 480826 362454
rect 481062 362218 481146 362454
rect 481382 362218 520826 362454
rect 521062 362218 521146 362454
rect 521382 362218 560826 362454
rect 561062 362218 561146 362454
rect 561382 362218 585342 362454
rect 585578 362218 585662 362454
rect 585898 362218 586890 362454
rect -2966 362134 586890 362218
rect -2966 361898 -1974 362134
rect -1738 361898 -1654 362134
rect -1418 361898 826 362134
rect 1062 361898 1146 362134
rect 1382 361898 40826 362134
rect 41062 361898 41146 362134
rect 41382 361898 80826 362134
rect 81062 361898 81146 362134
rect 81382 361898 120826 362134
rect 121062 361898 121146 362134
rect 121382 361898 160826 362134
rect 161062 361898 161146 362134
rect 161382 361898 200826 362134
rect 201062 361898 201146 362134
rect 201382 361898 240826 362134
rect 241062 361898 241146 362134
rect 241382 361898 280826 362134
rect 281062 361898 281146 362134
rect 281382 361898 320826 362134
rect 321062 361898 321146 362134
rect 321382 361898 360826 362134
rect 361062 361898 361146 362134
rect 361382 361898 400826 362134
rect 401062 361898 401146 362134
rect 401382 361898 440826 362134
rect 441062 361898 441146 362134
rect 441382 361898 480826 362134
rect 481062 361898 481146 362134
rect 481382 361898 520826 362134
rect 521062 361898 521146 362134
rect 521382 361898 560826 362134
rect 561062 361898 561146 362134
rect 561382 361898 585342 362134
rect 585578 361898 585662 362134
rect 585898 361898 586890 362134
rect -2966 361866 586890 361898
rect -8726 353614 592650 353646
rect -8726 353378 -8694 353614
rect -8458 353378 -8374 353614
rect -8138 353378 31986 353614
rect 32222 353378 32306 353614
rect 32542 353378 71986 353614
rect 72222 353378 72306 353614
rect 72542 353378 111986 353614
rect 112222 353378 112306 353614
rect 112542 353378 151986 353614
rect 152222 353378 152306 353614
rect 152542 353378 191986 353614
rect 192222 353378 192306 353614
rect 192542 353378 231986 353614
rect 232222 353378 232306 353614
rect 232542 353378 271986 353614
rect 272222 353378 272306 353614
rect 272542 353378 311986 353614
rect 312222 353378 312306 353614
rect 312542 353378 351986 353614
rect 352222 353378 352306 353614
rect 352542 353378 391986 353614
rect 392222 353378 392306 353614
rect 392542 353378 431986 353614
rect 432222 353378 432306 353614
rect 432542 353378 471986 353614
rect 472222 353378 472306 353614
rect 472542 353378 511986 353614
rect 512222 353378 512306 353614
rect 512542 353378 551986 353614
rect 552222 353378 552306 353614
rect 552542 353378 592062 353614
rect 592298 353378 592382 353614
rect 592618 353378 592650 353614
rect -8726 353294 592650 353378
rect -8726 353058 -8694 353294
rect -8458 353058 -8374 353294
rect -8138 353058 31986 353294
rect 32222 353058 32306 353294
rect 32542 353058 71986 353294
rect 72222 353058 72306 353294
rect 72542 353058 111986 353294
rect 112222 353058 112306 353294
rect 112542 353058 151986 353294
rect 152222 353058 152306 353294
rect 152542 353058 191986 353294
rect 192222 353058 192306 353294
rect 192542 353058 231986 353294
rect 232222 353058 232306 353294
rect 232542 353058 271986 353294
rect 272222 353058 272306 353294
rect 272542 353058 311986 353294
rect 312222 353058 312306 353294
rect 312542 353058 351986 353294
rect 352222 353058 352306 353294
rect 352542 353058 391986 353294
rect 392222 353058 392306 353294
rect 392542 353058 431986 353294
rect 432222 353058 432306 353294
rect 432542 353058 471986 353294
rect 472222 353058 472306 353294
rect 472542 353058 511986 353294
rect 512222 353058 512306 353294
rect 512542 353058 551986 353294
rect 552222 353058 552306 353294
rect 552542 353058 592062 353294
rect 592298 353058 592382 353294
rect 592618 353058 592650 353294
rect -8726 353026 592650 353058
rect -6806 349894 590730 349926
rect -6806 349658 -6774 349894
rect -6538 349658 -6454 349894
rect -6218 349658 28266 349894
rect 28502 349658 28586 349894
rect 28822 349658 68266 349894
rect 68502 349658 68586 349894
rect 68822 349658 108266 349894
rect 108502 349658 108586 349894
rect 108822 349658 148266 349894
rect 148502 349658 148586 349894
rect 148822 349658 188266 349894
rect 188502 349658 188586 349894
rect 188822 349658 228266 349894
rect 228502 349658 228586 349894
rect 228822 349658 268266 349894
rect 268502 349658 268586 349894
rect 268822 349658 308266 349894
rect 308502 349658 308586 349894
rect 308822 349658 348266 349894
rect 348502 349658 348586 349894
rect 348822 349658 388266 349894
rect 388502 349658 388586 349894
rect 388822 349658 428266 349894
rect 428502 349658 428586 349894
rect 428822 349658 468266 349894
rect 468502 349658 468586 349894
rect 468822 349658 508266 349894
rect 508502 349658 508586 349894
rect 508822 349658 548266 349894
rect 548502 349658 548586 349894
rect 548822 349658 590142 349894
rect 590378 349658 590462 349894
rect 590698 349658 590730 349894
rect -6806 349574 590730 349658
rect -6806 349338 -6774 349574
rect -6538 349338 -6454 349574
rect -6218 349338 28266 349574
rect 28502 349338 28586 349574
rect 28822 349338 68266 349574
rect 68502 349338 68586 349574
rect 68822 349338 108266 349574
rect 108502 349338 108586 349574
rect 108822 349338 148266 349574
rect 148502 349338 148586 349574
rect 148822 349338 188266 349574
rect 188502 349338 188586 349574
rect 188822 349338 228266 349574
rect 228502 349338 228586 349574
rect 228822 349338 268266 349574
rect 268502 349338 268586 349574
rect 268822 349338 308266 349574
rect 308502 349338 308586 349574
rect 308822 349338 348266 349574
rect 348502 349338 348586 349574
rect 348822 349338 388266 349574
rect 388502 349338 388586 349574
rect 388822 349338 428266 349574
rect 428502 349338 428586 349574
rect 428822 349338 468266 349574
rect 468502 349338 468586 349574
rect 468822 349338 508266 349574
rect 508502 349338 508586 349574
rect 508822 349338 548266 349574
rect 548502 349338 548586 349574
rect 548822 349338 590142 349574
rect 590378 349338 590462 349574
rect 590698 349338 590730 349574
rect -6806 349306 590730 349338
rect -4886 346174 588810 346206
rect -4886 345938 -4854 346174
rect -4618 345938 -4534 346174
rect -4298 345938 24546 346174
rect 24782 345938 24866 346174
rect 25102 345938 64546 346174
rect 64782 345938 64866 346174
rect 65102 345938 104546 346174
rect 104782 345938 104866 346174
rect 105102 345938 144546 346174
rect 144782 345938 144866 346174
rect 145102 345938 184546 346174
rect 184782 345938 184866 346174
rect 185102 345938 224546 346174
rect 224782 345938 224866 346174
rect 225102 345938 264546 346174
rect 264782 345938 264866 346174
rect 265102 345938 304546 346174
rect 304782 345938 304866 346174
rect 305102 345938 344546 346174
rect 344782 345938 344866 346174
rect 345102 345938 384546 346174
rect 384782 345938 384866 346174
rect 385102 345938 424546 346174
rect 424782 345938 424866 346174
rect 425102 345938 464546 346174
rect 464782 345938 464866 346174
rect 465102 345938 504546 346174
rect 504782 345938 504866 346174
rect 505102 345938 544546 346174
rect 544782 345938 544866 346174
rect 545102 345938 588222 346174
rect 588458 345938 588542 346174
rect 588778 345938 588810 346174
rect -4886 345854 588810 345938
rect -4886 345618 -4854 345854
rect -4618 345618 -4534 345854
rect -4298 345618 24546 345854
rect 24782 345618 24866 345854
rect 25102 345618 64546 345854
rect 64782 345618 64866 345854
rect 65102 345618 104546 345854
rect 104782 345618 104866 345854
rect 105102 345618 144546 345854
rect 144782 345618 144866 345854
rect 145102 345618 184546 345854
rect 184782 345618 184866 345854
rect 185102 345618 224546 345854
rect 224782 345618 224866 345854
rect 225102 345618 264546 345854
rect 264782 345618 264866 345854
rect 265102 345618 304546 345854
rect 304782 345618 304866 345854
rect 305102 345618 344546 345854
rect 344782 345618 344866 345854
rect 345102 345618 384546 345854
rect 384782 345618 384866 345854
rect 385102 345618 424546 345854
rect 424782 345618 424866 345854
rect 425102 345618 464546 345854
rect 464782 345618 464866 345854
rect 465102 345618 504546 345854
rect 504782 345618 504866 345854
rect 505102 345618 544546 345854
rect 544782 345618 544866 345854
rect 545102 345618 588222 345854
rect 588458 345618 588542 345854
rect 588778 345618 588810 345854
rect -4886 345586 588810 345618
rect -2966 342454 586890 342486
rect -2966 342218 -2934 342454
rect -2698 342218 -2614 342454
rect -2378 342218 20826 342454
rect 21062 342218 21146 342454
rect 21382 342218 60826 342454
rect 61062 342218 61146 342454
rect 61382 342218 100826 342454
rect 101062 342218 101146 342454
rect 101382 342218 140826 342454
rect 141062 342218 141146 342454
rect 141382 342218 180826 342454
rect 181062 342218 181146 342454
rect 181382 342218 220826 342454
rect 221062 342218 221146 342454
rect 221382 342218 260826 342454
rect 261062 342218 261146 342454
rect 261382 342218 300826 342454
rect 301062 342218 301146 342454
rect 301382 342218 340826 342454
rect 341062 342218 341146 342454
rect 341382 342218 380826 342454
rect 381062 342218 381146 342454
rect 381382 342218 420826 342454
rect 421062 342218 421146 342454
rect 421382 342218 460826 342454
rect 461062 342218 461146 342454
rect 461382 342218 500826 342454
rect 501062 342218 501146 342454
rect 501382 342218 540826 342454
rect 541062 342218 541146 342454
rect 541382 342218 580826 342454
rect 581062 342218 581146 342454
rect 581382 342218 586302 342454
rect 586538 342218 586622 342454
rect 586858 342218 586890 342454
rect -2966 342134 586890 342218
rect -2966 341898 -2934 342134
rect -2698 341898 -2614 342134
rect -2378 341898 20826 342134
rect 21062 341898 21146 342134
rect 21382 341898 60826 342134
rect 61062 341898 61146 342134
rect 61382 341898 100826 342134
rect 101062 341898 101146 342134
rect 101382 341898 140826 342134
rect 141062 341898 141146 342134
rect 141382 341898 180826 342134
rect 181062 341898 181146 342134
rect 181382 341898 220826 342134
rect 221062 341898 221146 342134
rect 221382 341898 260826 342134
rect 261062 341898 261146 342134
rect 261382 341898 300826 342134
rect 301062 341898 301146 342134
rect 301382 341898 340826 342134
rect 341062 341898 341146 342134
rect 341382 341898 380826 342134
rect 381062 341898 381146 342134
rect 381382 341898 420826 342134
rect 421062 341898 421146 342134
rect 421382 341898 460826 342134
rect 461062 341898 461146 342134
rect 461382 341898 500826 342134
rect 501062 341898 501146 342134
rect 501382 341898 540826 342134
rect 541062 341898 541146 342134
rect 541382 341898 580826 342134
rect 581062 341898 581146 342134
rect 581382 341898 586302 342134
rect 586538 341898 586622 342134
rect 586858 341898 586890 342134
rect -2966 341866 586890 341898
rect -8726 333614 592650 333646
rect -8726 333378 -7734 333614
rect -7498 333378 -7414 333614
rect -7178 333378 11986 333614
rect 12222 333378 12306 333614
rect 12542 333378 51986 333614
rect 52222 333378 52306 333614
rect 52542 333378 91986 333614
rect 92222 333378 92306 333614
rect 92542 333378 131986 333614
rect 132222 333378 132306 333614
rect 132542 333378 171986 333614
rect 172222 333378 172306 333614
rect 172542 333378 211986 333614
rect 212222 333378 212306 333614
rect 212542 333378 251986 333614
rect 252222 333378 252306 333614
rect 252542 333378 291986 333614
rect 292222 333378 292306 333614
rect 292542 333378 331986 333614
rect 332222 333378 332306 333614
rect 332542 333378 371986 333614
rect 372222 333378 372306 333614
rect 372542 333378 411986 333614
rect 412222 333378 412306 333614
rect 412542 333378 451986 333614
rect 452222 333378 452306 333614
rect 452542 333378 491986 333614
rect 492222 333378 492306 333614
rect 492542 333378 531986 333614
rect 532222 333378 532306 333614
rect 532542 333378 571986 333614
rect 572222 333378 572306 333614
rect 572542 333378 591102 333614
rect 591338 333378 591422 333614
rect 591658 333378 592650 333614
rect -8726 333294 592650 333378
rect -8726 333058 -7734 333294
rect -7498 333058 -7414 333294
rect -7178 333058 11986 333294
rect 12222 333058 12306 333294
rect 12542 333058 51986 333294
rect 52222 333058 52306 333294
rect 52542 333058 91986 333294
rect 92222 333058 92306 333294
rect 92542 333058 131986 333294
rect 132222 333058 132306 333294
rect 132542 333058 171986 333294
rect 172222 333058 172306 333294
rect 172542 333058 211986 333294
rect 212222 333058 212306 333294
rect 212542 333058 251986 333294
rect 252222 333058 252306 333294
rect 252542 333058 291986 333294
rect 292222 333058 292306 333294
rect 292542 333058 331986 333294
rect 332222 333058 332306 333294
rect 332542 333058 371986 333294
rect 372222 333058 372306 333294
rect 372542 333058 411986 333294
rect 412222 333058 412306 333294
rect 412542 333058 451986 333294
rect 452222 333058 452306 333294
rect 452542 333058 491986 333294
rect 492222 333058 492306 333294
rect 492542 333058 531986 333294
rect 532222 333058 532306 333294
rect 532542 333058 571986 333294
rect 572222 333058 572306 333294
rect 572542 333058 591102 333294
rect 591338 333058 591422 333294
rect 591658 333058 592650 333294
rect -8726 333026 592650 333058
rect -6806 329894 590730 329926
rect -6806 329658 -5814 329894
rect -5578 329658 -5494 329894
rect -5258 329658 8266 329894
rect 8502 329658 8586 329894
rect 8822 329658 48266 329894
rect 48502 329658 48586 329894
rect 48822 329658 88266 329894
rect 88502 329658 88586 329894
rect 88822 329658 128266 329894
rect 128502 329658 128586 329894
rect 128822 329658 168266 329894
rect 168502 329658 168586 329894
rect 168822 329658 208266 329894
rect 208502 329658 208586 329894
rect 208822 329658 248266 329894
rect 248502 329658 248586 329894
rect 248822 329658 288266 329894
rect 288502 329658 288586 329894
rect 288822 329658 328266 329894
rect 328502 329658 328586 329894
rect 328822 329658 368266 329894
rect 368502 329658 368586 329894
rect 368822 329658 408266 329894
rect 408502 329658 408586 329894
rect 408822 329658 448266 329894
rect 448502 329658 448586 329894
rect 448822 329658 488266 329894
rect 488502 329658 488586 329894
rect 488822 329658 528266 329894
rect 528502 329658 528586 329894
rect 528822 329658 568266 329894
rect 568502 329658 568586 329894
rect 568822 329658 589182 329894
rect 589418 329658 589502 329894
rect 589738 329658 590730 329894
rect -6806 329574 590730 329658
rect -6806 329338 -5814 329574
rect -5578 329338 -5494 329574
rect -5258 329338 8266 329574
rect 8502 329338 8586 329574
rect 8822 329338 48266 329574
rect 48502 329338 48586 329574
rect 48822 329338 88266 329574
rect 88502 329338 88586 329574
rect 88822 329338 128266 329574
rect 128502 329338 128586 329574
rect 128822 329338 168266 329574
rect 168502 329338 168586 329574
rect 168822 329338 208266 329574
rect 208502 329338 208586 329574
rect 208822 329338 248266 329574
rect 248502 329338 248586 329574
rect 248822 329338 288266 329574
rect 288502 329338 288586 329574
rect 288822 329338 328266 329574
rect 328502 329338 328586 329574
rect 328822 329338 368266 329574
rect 368502 329338 368586 329574
rect 368822 329338 408266 329574
rect 408502 329338 408586 329574
rect 408822 329338 448266 329574
rect 448502 329338 448586 329574
rect 448822 329338 488266 329574
rect 488502 329338 488586 329574
rect 488822 329338 528266 329574
rect 528502 329338 528586 329574
rect 528822 329338 568266 329574
rect 568502 329338 568586 329574
rect 568822 329338 589182 329574
rect 589418 329338 589502 329574
rect 589738 329338 590730 329574
rect -6806 329306 590730 329338
rect -4886 326174 588810 326206
rect -4886 325938 -3894 326174
rect -3658 325938 -3574 326174
rect -3338 325938 4546 326174
rect 4782 325938 4866 326174
rect 5102 325938 44546 326174
rect 44782 325938 44866 326174
rect 45102 325938 84546 326174
rect 84782 325938 84866 326174
rect 85102 325938 124546 326174
rect 124782 325938 124866 326174
rect 125102 325938 164546 326174
rect 164782 325938 164866 326174
rect 165102 325938 204546 326174
rect 204782 325938 204866 326174
rect 205102 325938 244546 326174
rect 244782 325938 244866 326174
rect 245102 325938 284546 326174
rect 284782 325938 284866 326174
rect 285102 325938 324546 326174
rect 324782 325938 324866 326174
rect 325102 325938 364546 326174
rect 364782 325938 364866 326174
rect 365102 325938 404546 326174
rect 404782 325938 404866 326174
rect 405102 325938 444546 326174
rect 444782 325938 444866 326174
rect 445102 325938 484546 326174
rect 484782 325938 484866 326174
rect 485102 325938 524546 326174
rect 524782 325938 524866 326174
rect 525102 325938 564546 326174
rect 564782 325938 564866 326174
rect 565102 325938 587262 326174
rect 587498 325938 587582 326174
rect 587818 325938 588810 326174
rect -4886 325854 588810 325938
rect -4886 325618 -3894 325854
rect -3658 325618 -3574 325854
rect -3338 325618 4546 325854
rect 4782 325618 4866 325854
rect 5102 325618 44546 325854
rect 44782 325618 44866 325854
rect 45102 325618 84546 325854
rect 84782 325618 84866 325854
rect 85102 325618 124546 325854
rect 124782 325618 124866 325854
rect 125102 325618 164546 325854
rect 164782 325618 164866 325854
rect 165102 325618 204546 325854
rect 204782 325618 204866 325854
rect 205102 325618 244546 325854
rect 244782 325618 244866 325854
rect 245102 325618 284546 325854
rect 284782 325618 284866 325854
rect 285102 325618 324546 325854
rect 324782 325618 324866 325854
rect 325102 325618 364546 325854
rect 364782 325618 364866 325854
rect 365102 325618 404546 325854
rect 404782 325618 404866 325854
rect 405102 325618 444546 325854
rect 444782 325618 444866 325854
rect 445102 325618 484546 325854
rect 484782 325618 484866 325854
rect 485102 325618 524546 325854
rect 524782 325618 524866 325854
rect 525102 325618 564546 325854
rect 564782 325618 564866 325854
rect 565102 325618 587262 325854
rect 587498 325618 587582 325854
rect 587818 325618 588810 325854
rect -4886 325586 588810 325618
rect -2966 322454 586890 322486
rect -2966 322218 -1974 322454
rect -1738 322218 -1654 322454
rect -1418 322218 826 322454
rect 1062 322218 1146 322454
rect 1382 322218 40826 322454
rect 41062 322218 41146 322454
rect 41382 322218 80826 322454
rect 81062 322218 81146 322454
rect 81382 322218 120826 322454
rect 121062 322218 121146 322454
rect 121382 322218 160826 322454
rect 161062 322218 161146 322454
rect 161382 322218 200826 322454
rect 201062 322218 201146 322454
rect 201382 322218 240826 322454
rect 241062 322218 241146 322454
rect 241382 322218 280826 322454
rect 281062 322218 281146 322454
rect 281382 322218 320826 322454
rect 321062 322218 321146 322454
rect 321382 322218 360826 322454
rect 361062 322218 361146 322454
rect 361382 322218 400826 322454
rect 401062 322218 401146 322454
rect 401382 322218 440826 322454
rect 441062 322218 441146 322454
rect 441382 322218 480826 322454
rect 481062 322218 481146 322454
rect 481382 322218 520826 322454
rect 521062 322218 521146 322454
rect 521382 322218 560826 322454
rect 561062 322218 561146 322454
rect 561382 322218 585342 322454
rect 585578 322218 585662 322454
rect 585898 322218 586890 322454
rect -2966 322134 586890 322218
rect -2966 321898 -1974 322134
rect -1738 321898 -1654 322134
rect -1418 321898 826 322134
rect 1062 321898 1146 322134
rect 1382 321898 40826 322134
rect 41062 321898 41146 322134
rect 41382 321898 80826 322134
rect 81062 321898 81146 322134
rect 81382 321898 120826 322134
rect 121062 321898 121146 322134
rect 121382 321898 160826 322134
rect 161062 321898 161146 322134
rect 161382 321898 200826 322134
rect 201062 321898 201146 322134
rect 201382 321898 240826 322134
rect 241062 321898 241146 322134
rect 241382 321898 280826 322134
rect 281062 321898 281146 322134
rect 281382 321898 320826 322134
rect 321062 321898 321146 322134
rect 321382 321898 360826 322134
rect 361062 321898 361146 322134
rect 361382 321898 400826 322134
rect 401062 321898 401146 322134
rect 401382 321898 440826 322134
rect 441062 321898 441146 322134
rect 441382 321898 480826 322134
rect 481062 321898 481146 322134
rect 481382 321898 520826 322134
rect 521062 321898 521146 322134
rect 521382 321898 560826 322134
rect 561062 321898 561146 322134
rect 561382 321898 585342 322134
rect 585578 321898 585662 322134
rect 585898 321898 586890 322134
rect -2966 321866 586890 321898
rect -8726 313614 592650 313646
rect -8726 313378 -8694 313614
rect -8458 313378 -8374 313614
rect -8138 313378 31986 313614
rect 32222 313378 32306 313614
rect 32542 313378 71986 313614
rect 72222 313378 72306 313614
rect 72542 313378 111986 313614
rect 112222 313378 112306 313614
rect 112542 313378 151986 313614
rect 152222 313378 152306 313614
rect 152542 313378 191986 313614
rect 192222 313378 192306 313614
rect 192542 313378 231986 313614
rect 232222 313378 232306 313614
rect 232542 313378 271986 313614
rect 272222 313378 272306 313614
rect 272542 313378 311986 313614
rect 312222 313378 312306 313614
rect 312542 313378 351986 313614
rect 352222 313378 352306 313614
rect 352542 313378 391986 313614
rect 392222 313378 392306 313614
rect 392542 313378 431986 313614
rect 432222 313378 432306 313614
rect 432542 313378 471986 313614
rect 472222 313378 472306 313614
rect 472542 313378 511986 313614
rect 512222 313378 512306 313614
rect 512542 313378 551986 313614
rect 552222 313378 552306 313614
rect 552542 313378 592062 313614
rect 592298 313378 592382 313614
rect 592618 313378 592650 313614
rect -8726 313294 592650 313378
rect -8726 313058 -8694 313294
rect -8458 313058 -8374 313294
rect -8138 313058 31986 313294
rect 32222 313058 32306 313294
rect 32542 313058 71986 313294
rect 72222 313058 72306 313294
rect 72542 313058 111986 313294
rect 112222 313058 112306 313294
rect 112542 313058 151986 313294
rect 152222 313058 152306 313294
rect 152542 313058 191986 313294
rect 192222 313058 192306 313294
rect 192542 313058 231986 313294
rect 232222 313058 232306 313294
rect 232542 313058 271986 313294
rect 272222 313058 272306 313294
rect 272542 313058 311986 313294
rect 312222 313058 312306 313294
rect 312542 313058 351986 313294
rect 352222 313058 352306 313294
rect 352542 313058 391986 313294
rect 392222 313058 392306 313294
rect 392542 313058 431986 313294
rect 432222 313058 432306 313294
rect 432542 313058 471986 313294
rect 472222 313058 472306 313294
rect 472542 313058 511986 313294
rect 512222 313058 512306 313294
rect 512542 313058 551986 313294
rect 552222 313058 552306 313294
rect 552542 313058 592062 313294
rect 592298 313058 592382 313294
rect 592618 313058 592650 313294
rect -8726 313026 592650 313058
rect -6806 309894 590730 309926
rect -6806 309658 -6774 309894
rect -6538 309658 -6454 309894
rect -6218 309658 28266 309894
rect 28502 309658 28586 309894
rect 28822 309658 68266 309894
rect 68502 309658 68586 309894
rect 68822 309658 108266 309894
rect 108502 309658 108586 309894
rect 108822 309658 148266 309894
rect 148502 309658 148586 309894
rect 148822 309658 188266 309894
rect 188502 309658 188586 309894
rect 188822 309658 228266 309894
rect 228502 309658 228586 309894
rect 228822 309658 268266 309894
rect 268502 309658 268586 309894
rect 268822 309658 308266 309894
rect 308502 309658 308586 309894
rect 308822 309658 348266 309894
rect 348502 309658 348586 309894
rect 348822 309658 388266 309894
rect 388502 309658 388586 309894
rect 388822 309658 428266 309894
rect 428502 309658 428586 309894
rect 428822 309658 468266 309894
rect 468502 309658 468586 309894
rect 468822 309658 508266 309894
rect 508502 309658 508586 309894
rect 508822 309658 548266 309894
rect 548502 309658 548586 309894
rect 548822 309658 590142 309894
rect 590378 309658 590462 309894
rect 590698 309658 590730 309894
rect -6806 309574 590730 309658
rect -6806 309338 -6774 309574
rect -6538 309338 -6454 309574
rect -6218 309338 28266 309574
rect 28502 309338 28586 309574
rect 28822 309338 68266 309574
rect 68502 309338 68586 309574
rect 68822 309338 108266 309574
rect 108502 309338 108586 309574
rect 108822 309338 148266 309574
rect 148502 309338 148586 309574
rect 148822 309338 188266 309574
rect 188502 309338 188586 309574
rect 188822 309338 228266 309574
rect 228502 309338 228586 309574
rect 228822 309338 268266 309574
rect 268502 309338 268586 309574
rect 268822 309338 308266 309574
rect 308502 309338 308586 309574
rect 308822 309338 348266 309574
rect 348502 309338 348586 309574
rect 348822 309338 388266 309574
rect 388502 309338 388586 309574
rect 388822 309338 428266 309574
rect 428502 309338 428586 309574
rect 428822 309338 468266 309574
rect 468502 309338 468586 309574
rect 468822 309338 508266 309574
rect 508502 309338 508586 309574
rect 508822 309338 548266 309574
rect 548502 309338 548586 309574
rect 548822 309338 590142 309574
rect 590378 309338 590462 309574
rect 590698 309338 590730 309574
rect -6806 309306 590730 309338
rect -4886 306174 588810 306206
rect -4886 305938 -4854 306174
rect -4618 305938 -4534 306174
rect -4298 305938 24546 306174
rect 24782 305938 24866 306174
rect 25102 305938 64546 306174
rect 64782 305938 64866 306174
rect 65102 305938 104546 306174
rect 104782 305938 104866 306174
rect 105102 305938 144546 306174
rect 144782 305938 144866 306174
rect 145102 305938 184546 306174
rect 184782 305938 184866 306174
rect 185102 305938 224546 306174
rect 224782 305938 224866 306174
rect 225102 305938 264546 306174
rect 264782 305938 264866 306174
rect 265102 305938 304546 306174
rect 304782 305938 304866 306174
rect 305102 305938 344546 306174
rect 344782 305938 344866 306174
rect 345102 305938 384546 306174
rect 384782 305938 384866 306174
rect 385102 305938 424546 306174
rect 424782 305938 424866 306174
rect 425102 305938 464546 306174
rect 464782 305938 464866 306174
rect 465102 305938 504546 306174
rect 504782 305938 504866 306174
rect 505102 305938 544546 306174
rect 544782 305938 544866 306174
rect 545102 305938 588222 306174
rect 588458 305938 588542 306174
rect 588778 305938 588810 306174
rect -4886 305854 588810 305938
rect -4886 305618 -4854 305854
rect -4618 305618 -4534 305854
rect -4298 305618 24546 305854
rect 24782 305618 24866 305854
rect 25102 305618 64546 305854
rect 64782 305618 64866 305854
rect 65102 305618 104546 305854
rect 104782 305618 104866 305854
rect 105102 305618 144546 305854
rect 144782 305618 144866 305854
rect 145102 305618 184546 305854
rect 184782 305618 184866 305854
rect 185102 305618 224546 305854
rect 224782 305618 224866 305854
rect 225102 305618 264546 305854
rect 264782 305618 264866 305854
rect 265102 305618 304546 305854
rect 304782 305618 304866 305854
rect 305102 305618 344546 305854
rect 344782 305618 344866 305854
rect 345102 305618 384546 305854
rect 384782 305618 384866 305854
rect 385102 305618 424546 305854
rect 424782 305618 424866 305854
rect 425102 305618 464546 305854
rect 464782 305618 464866 305854
rect 465102 305618 504546 305854
rect 504782 305618 504866 305854
rect 505102 305618 544546 305854
rect 544782 305618 544866 305854
rect 545102 305618 588222 305854
rect 588458 305618 588542 305854
rect 588778 305618 588810 305854
rect -4886 305586 588810 305618
rect -2966 302454 586890 302486
rect -2966 302218 -2934 302454
rect -2698 302218 -2614 302454
rect -2378 302218 20826 302454
rect 21062 302218 21146 302454
rect 21382 302218 60826 302454
rect 61062 302218 61146 302454
rect 61382 302218 100826 302454
rect 101062 302218 101146 302454
rect 101382 302218 140826 302454
rect 141382 302218 180826 302454
rect 181382 302218 220826 302454
rect 221382 302218 260826 302454
rect 261382 302218 300826 302454
rect 301382 302218 340826 302454
rect 341062 302218 341146 302454
rect 341382 302218 380826 302454
rect 381062 302218 381146 302454
rect 381382 302218 420826 302454
rect 421062 302218 421146 302454
rect 421382 302218 460826 302454
rect 461062 302218 461146 302454
rect 461382 302218 500826 302454
rect 501062 302218 501146 302454
rect 501382 302218 540826 302454
rect 541062 302218 541146 302454
rect 541382 302218 580826 302454
rect 581062 302218 581146 302454
rect 581382 302218 586302 302454
rect 586538 302218 586622 302454
rect 586858 302218 586890 302454
rect -2966 302134 586890 302218
rect -2966 301898 -2934 302134
rect -2698 301898 -2614 302134
rect -2378 301898 20826 302134
rect 21062 301898 21146 302134
rect 21382 301898 60826 302134
rect 61062 301898 61146 302134
rect 61382 301898 100826 302134
rect 101062 301898 101146 302134
rect 101382 301898 140826 302134
rect 141382 301898 180826 302134
rect 181382 301898 220826 302134
rect 221382 301898 260826 302134
rect 261382 301898 300826 302134
rect 301382 301898 340826 302134
rect 341062 301898 341146 302134
rect 341382 301898 380826 302134
rect 381062 301898 381146 302134
rect 381382 301898 420826 302134
rect 421062 301898 421146 302134
rect 421382 301898 460826 302134
rect 461062 301898 461146 302134
rect 461382 301898 500826 302134
rect 501062 301898 501146 302134
rect 501382 301898 540826 302134
rect 541062 301898 541146 302134
rect 541382 301898 580826 302134
rect 581062 301898 581146 302134
rect 581382 301898 586302 302134
rect 586538 301898 586622 302134
rect 586858 301898 586890 302134
rect -2966 301866 586890 301898
rect -8726 293614 592650 293646
rect -8726 293378 -7734 293614
rect -7498 293378 -7414 293614
rect -7178 293378 11986 293614
rect 12222 293378 12306 293614
rect 12542 293378 51986 293614
rect 52222 293378 52306 293614
rect 52542 293378 91986 293614
rect 92222 293378 92306 293614
rect 92542 293378 131986 293614
rect 132222 293378 132306 293614
rect 132542 293378 171986 293614
rect 172222 293378 172306 293614
rect 172542 293378 211986 293614
rect 212222 293378 212306 293614
rect 212542 293378 251986 293614
rect 252222 293378 252306 293614
rect 252542 293378 291986 293614
rect 292222 293378 292306 293614
rect 292542 293378 331986 293614
rect 332222 293378 332306 293614
rect 332542 293378 371986 293614
rect 372222 293378 372306 293614
rect 372542 293378 411986 293614
rect 412222 293378 412306 293614
rect 412542 293378 451986 293614
rect 452222 293378 452306 293614
rect 452542 293378 491986 293614
rect 492222 293378 492306 293614
rect 492542 293378 531986 293614
rect 532222 293378 532306 293614
rect 532542 293378 571986 293614
rect 572222 293378 572306 293614
rect 572542 293378 591102 293614
rect 591338 293378 591422 293614
rect 591658 293378 592650 293614
rect -8726 293294 592650 293378
rect -8726 293058 -7734 293294
rect -7498 293058 -7414 293294
rect -7178 293058 11986 293294
rect 12222 293058 12306 293294
rect 12542 293058 51986 293294
rect 52222 293058 52306 293294
rect 52542 293058 91986 293294
rect 92222 293058 92306 293294
rect 92542 293058 131986 293294
rect 132222 293058 132306 293294
rect 132542 293058 171986 293294
rect 172222 293058 172306 293294
rect 172542 293058 211986 293294
rect 212222 293058 212306 293294
rect 212542 293058 251986 293294
rect 252222 293058 252306 293294
rect 252542 293058 291986 293294
rect 292222 293058 292306 293294
rect 292542 293058 331986 293294
rect 332222 293058 332306 293294
rect 332542 293058 371986 293294
rect 372222 293058 372306 293294
rect 372542 293058 411986 293294
rect 412222 293058 412306 293294
rect 412542 293058 451986 293294
rect 452222 293058 452306 293294
rect 452542 293058 491986 293294
rect 492222 293058 492306 293294
rect 492542 293058 531986 293294
rect 532222 293058 532306 293294
rect 532542 293058 571986 293294
rect 572222 293058 572306 293294
rect 572542 293058 591102 293294
rect 591338 293058 591422 293294
rect 591658 293058 592650 293294
rect -8726 293026 592650 293058
rect -6806 289894 590730 289926
rect -6806 289658 -5814 289894
rect -5578 289658 -5494 289894
rect -5258 289658 8266 289894
rect 8502 289658 8586 289894
rect 8822 289658 48266 289894
rect 48502 289658 48586 289894
rect 48822 289658 88266 289894
rect 88502 289658 88586 289894
rect 88822 289658 128266 289894
rect 128502 289658 128586 289894
rect 128822 289658 168266 289894
rect 168502 289658 168586 289894
rect 168822 289658 208266 289894
rect 208502 289658 208586 289894
rect 208822 289658 248266 289894
rect 248502 289658 248586 289894
rect 248822 289658 288266 289894
rect 288502 289658 288586 289894
rect 288822 289658 328266 289894
rect 328502 289658 328586 289894
rect 328822 289658 368266 289894
rect 368502 289658 368586 289894
rect 368822 289658 408266 289894
rect 408502 289658 408586 289894
rect 408822 289658 448266 289894
rect 448502 289658 448586 289894
rect 448822 289658 488266 289894
rect 488502 289658 488586 289894
rect 488822 289658 528266 289894
rect 528502 289658 528586 289894
rect 528822 289658 568266 289894
rect 568502 289658 568586 289894
rect 568822 289658 589182 289894
rect 589418 289658 589502 289894
rect 589738 289658 590730 289894
rect -6806 289574 590730 289658
rect -6806 289338 -5814 289574
rect -5578 289338 -5494 289574
rect -5258 289338 8266 289574
rect 8502 289338 8586 289574
rect 8822 289338 48266 289574
rect 48502 289338 48586 289574
rect 48822 289338 88266 289574
rect 88502 289338 88586 289574
rect 88822 289338 128266 289574
rect 128502 289338 128586 289574
rect 128822 289338 168266 289574
rect 168502 289338 168586 289574
rect 168822 289338 208266 289574
rect 208502 289338 208586 289574
rect 208822 289338 248266 289574
rect 248502 289338 248586 289574
rect 248822 289338 288266 289574
rect 288502 289338 288586 289574
rect 288822 289338 328266 289574
rect 328502 289338 328586 289574
rect 328822 289338 368266 289574
rect 368502 289338 368586 289574
rect 368822 289338 408266 289574
rect 408502 289338 408586 289574
rect 408822 289338 448266 289574
rect 448502 289338 448586 289574
rect 448822 289338 488266 289574
rect 488502 289338 488586 289574
rect 488822 289338 528266 289574
rect 528502 289338 528586 289574
rect 528822 289338 568266 289574
rect 568502 289338 568586 289574
rect 568822 289338 589182 289574
rect 589418 289338 589502 289574
rect 589738 289338 590730 289574
rect -6806 289306 590730 289338
rect -4886 286174 588810 286206
rect -4886 285938 -3894 286174
rect -3658 285938 -3574 286174
rect -3338 285938 4546 286174
rect 4782 285938 4866 286174
rect 5102 285938 44546 286174
rect 44782 285938 44866 286174
rect 45102 285938 84546 286174
rect 84782 285938 84866 286174
rect 85102 285938 124546 286174
rect 124782 285938 124866 286174
rect 125102 285938 164546 286174
rect 164782 285938 164866 286174
rect 165102 285938 204546 286174
rect 204782 285938 204866 286174
rect 205102 285938 244546 286174
rect 244782 285938 244866 286174
rect 245102 285938 284546 286174
rect 284782 285938 284866 286174
rect 285102 285938 324546 286174
rect 324782 285938 324866 286174
rect 325102 285938 364546 286174
rect 364782 285938 364866 286174
rect 365102 285938 404546 286174
rect 404782 285938 404866 286174
rect 405102 285938 444546 286174
rect 444782 285938 444866 286174
rect 445102 285938 484546 286174
rect 484782 285938 484866 286174
rect 485102 285938 524546 286174
rect 524782 285938 524866 286174
rect 525102 285938 564546 286174
rect 564782 285938 564866 286174
rect 565102 285938 587262 286174
rect 587498 285938 587582 286174
rect 587818 285938 588810 286174
rect -4886 285854 588810 285938
rect -4886 285618 -3894 285854
rect -3658 285618 -3574 285854
rect -3338 285618 4546 285854
rect 4782 285618 4866 285854
rect 5102 285618 44546 285854
rect 44782 285618 44866 285854
rect 45102 285618 84546 285854
rect 84782 285618 84866 285854
rect 85102 285618 124546 285854
rect 124782 285618 124866 285854
rect 125102 285618 164546 285854
rect 164782 285618 164866 285854
rect 165102 285618 204546 285854
rect 204782 285618 204866 285854
rect 205102 285618 244546 285854
rect 244782 285618 244866 285854
rect 245102 285618 284546 285854
rect 284782 285618 284866 285854
rect 285102 285618 324546 285854
rect 324782 285618 324866 285854
rect 325102 285618 364546 285854
rect 364782 285618 364866 285854
rect 365102 285618 404546 285854
rect 404782 285618 404866 285854
rect 405102 285618 444546 285854
rect 444782 285618 444866 285854
rect 445102 285618 484546 285854
rect 484782 285618 484866 285854
rect 485102 285618 524546 285854
rect 524782 285618 524866 285854
rect 525102 285618 564546 285854
rect 564782 285618 564866 285854
rect 565102 285618 587262 285854
rect 587498 285618 587582 285854
rect 587818 285618 588810 285854
rect -4886 285586 588810 285618
rect -2966 282454 586890 282486
rect -2966 282218 -1974 282454
rect -1738 282218 -1654 282454
rect -1418 282218 826 282454
rect 1062 282218 1146 282454
rect 1382 282218 40826 282454
rect 41062 282218 41146 282454
rect 41382 282218 80826 282454
rect 81062 282218 81146 282454
rect 81382 282218 120826 282454
rect 121062 282218 121146 282454
rect 121382 282218 160826 282454
rect 161382 282218 200826 282454
rect 201382 282218 240826 282454
rect 241382 282218 280826 282454
rect 281382 282218 320826 282454
rect 321062 282218 321146 282454
rect 321382 282218 360826 282454
rect 361062 282218 361146 282454
rect 361382 282218 400826 282454
rect 401062 282218 401146 282454
rect 401382 282218 440826 282454
rect 441062 282218 441146 282454
rect 441382 282218 480826 282454
rect 481062 282218 481146 282454
rect 481382 282218 520826 282454
rect 521062 282218 521146 282454
rect 521382 282218 560826 282454
rect 561062 282218 561146 282454
rect 561382 282218 585342 282454
rect 585578 282218 585662 282454
rect 585898 282218 586890 282454
rect -2966 282134 586890 282218
rect -2966 281898 -1974 282134
rect -1738 281898 -1654 282134
rect -1418 281898 826 282134
rect 1062 281898 1146 282134
rect 1382 281898 40826 282134
rect 41062 281898 41146 282134
rect 41382 281898 80826 282134
rect 81062 281898 81146 282134
rect 81382 281898 120826 282134
rect 121062 281898 121146 282134
rect 121382 281898 160826 282134
rect 161382 281898 200826 282134
rect 201382 281898 240826 282134
rect 241382 281898 280826 282134
rect 281382 281898 320826 282134
rect 321062 281898 321146 282134
rect 321382 281898 360826 282134
rect 361062 281898 361146 282134
rect 361382 281898 400826 282134
rect 401062 281898 401146 282134
rect 401382 281898 440826 282134
rect 441062 281898 441146 282134
rect 441382 281898 480826 282134
rect 481062 281898 481146 282134
rect 481382 281898 520826 282134
rect 521062 281898 521146 282134
rect 521382 281898 560826 282134
rect 561062 281898 561146 282134
rect 561382 281898 585342 282134
rect 585578 281898 585662 282134
rect 585898 281898 586890 282134
rect -2966 281866 586890 281898
rect -8726 273614 592650 273646
rect -8726 273378 -8694 273614
rect -8458 273378 -8374 273614
rect -8138 273378 31986 273614
rect 32222 273378 32306 273614
rect 32542 273378 71986 273614
rect 72222 273378 72306 273614
rect 72542 273378 111986 273614
rect 112222 273378 112306 273614
rect 112542 273378 151986 273614
rect 152222 273378 152306 273614
rect 152542 273378 191986 273614
rect 192222 273378 192306 273614
rect 192542 273378 231986 273614
rect 232222 273378 232306 273614
rect 232542 273378 271986 273614
rect 272222 273378 272306 273614
rect 272542 273378 311986 273614
rect 312222 273378 312306 273614
rect 312542 273378 351986 273614
rect 352222 273378 352306 273614
rect 352542 273378 391986 273614
rect 392222 273378 392306 273614
rect 392542 273378 431986 273614
rect 432222 273378 432306 273614
rect 432542 273378 471986 273614
rect 472222 273378 472306 273614
rect 472542 273378 511986 273614
rect 512222 273378 512306 273614
rect 512542 273378 551986 273614
rect 552222 273378 552306 273614
rect 552542 273378 592062 273614
rect 592298 273378 592382 273614
rect 592618 273378 592650 273614
rect -8726 273294 592650 273378
rect -8726 273058 -8694 273294
rect -8458 273058 -8374 273294
rect -8138 273058 31986 273294
rect 32222 273058 32306 273294
rect 32542 273058 71986 273294
rect 72222 273058 72306 273294
rect 72542 273058 111986 273294
rect 112222 273058 112306 273294
rect 112542 273058 151986 273294
rect 152222 273058 152306 273294
rect 152542 273058 191986 273294
rect 192222 273058 192306 273294
rect 192542 273058 231986 273294
rect 232222 273058 232306 273294
rect 232542 273058 271986 273294
rect 272222 273058 272306 273294
rect 272542 273058 311986 273294
rect 312222 273058 312306 273294
rect 312542 273058 351986 273294
rect 352222 273058 352306 273294
rect 352542 273058 391986 273294
rect 392222 273058 392306 273294
rect 392542 273058 431986 273294
rect 432222 273058 432306 273294
rect 432542 273058 471986 273294
rect 472222 273058 472306 273294
rect 472542 273058 511986 273294
rect 512222 273058 512306 273294
rect 512542 273058 551986 273294
rect 552222 273058 552306 273294
rect 552542 273058 592062 273294
rect 592298 273058 592382 273294
rect 592618 273058 592650 273294
rect -8726 273026 592650 273058
rect -6806 269894 590730 269926
rect -6806 269658 -6774 269894
rect -6538 269658 -6454 269894
rect -6218 269658 28266 269894
rect 28502 269658 28586 269894
rect 28822 269658 68266 269894
rect 68502 269658 68586 269894
rect 68822 269658 108266 269894
rect 108502 269658 108586 269894
rect 108822 269658 148266 269894
rect 148502 269658 148586 269894
rect 148822 269658 188266 269894
rect 188502 269658 188586 269894
rect 188822 269658 228266 269894
rect 228502 269658 228586 269894
rect 228822 269658 268266 269894
rect 268502 269658 268586 269894
rect 268822 269658 308266 269894
rect 308502 269658 308586 269894
rect 308822 269658 348266 269894
rect 348502 269658 348586 269894
rect 348822 269658 388266 269894
rect 388502 269658 388586 269894
rect 388822 269658 428266 269894
rect 428502 269658 428586 269894
rect 428822 269658 468266 269894
rect 468502 269658 468586 269894
rect 468822 269658 508266 269894
rect 508502 269658 508586 269894
rect 508822 269658 548266 269894
rect 548502 269658 548586 269894
rect 548822 269658 590142 269894
rect 590378 269658 590462 269894
rect 590698 269658 590730 269894
rect -6806 269574 590730 269658
rect -6806 269338 -6774 269574
rect -6538 269338 -6454 269574
rect -6218 269338 28266 269574
rect 28502 269338 28586 269574
rect 28822 269338 68266 269574
rect 68502 269338 68586 269574
rect 68822 269338 108266 269574
rect 108502 269338 108586 269574
rect 108822 269338 148266 269574
rect 148502 269338 148586 269574
rect 148822 269338 188266 269574
rect 188502 269338 188586 269574
rect 188822 269338 228266 269574
rect 228502 269338 228586 269574
rect 228822 269338 268266 269574
rect 268502 269338 268586 269574
rect 268822 269338 308266 269574
rect 308502 269338 308586 269574
rect 308822 269338 348266 269574
rect 348502 269338 348586 269574
rect 348822 269338 388266 269574
rect 388502 269338 388586 269574
rect 388822 269338 428266 269574
rect 428502 269338 428586 269574
rect 428822 269338 468266 269574
rect 468502 269338 468586 269574
rect 468822 269338 508266 269574
rect 508502 269338 508586 269574
rect 508822 269338 548266 269574
rect 548502 269338 548586 269574
rect 548822 269338 590142 269574
rect 590378 269338 590462 269574
rect 590698 269338 590730 269574
rect -6806 269306 590730 269338
rect -4886 266174 588810 266206
rect -4886 265938 -4854 266174
rect -4618 265938 -4534 266174
rect -4298 265938 24546 266174
rect 24782 265938 24866 266174
rect 25102 265938 64546 266174
rect 64782 265938 64866 266174
rect 65102 265938 104546 266174
rect 104782 265938 104866 266174
rect 105102 265938 144546 266174
rect 144782 265938 144866 266174
rect 145102 265938 184546 266174
rect 184782 265938 184866 266174
rect 185102 265938 224546 266174
rect 224782 265938 224866 266174
rect 225102 265938 264546 266174
rect 264782 265938 264866 266174
rect 265102 265938 304546 266174
rect 304782 265938 304866 266174
rect 305102 265938 344546 266174
rect 344782 265938 344866 266174
rect 345102 265938 384546 266174
rect 384782 265938 384866 266174
rect 385102 265938 424546 266174
rect 424782 265938 424866 266174
rect 425102 265938 464546 266174
rect 464782 265938 464866 266174
rect 465102 265938 504546 266174
rect 504782 265938 504866 266174
rect 505102 265938 544546 266174
rect 544782 265938 544866 266174
rect 545102 265938 588222 266174
rect 588458 265938 588542 266174
rect 588778 265938 588810 266174
rect -4886 265854 588810 265938
rect -4886 265618 -4854 265854
rect -4618 265618 -4534 265854
rect -4298 265618 24546 265854
rect 24782 265618 24866 265854
rect 25102 265618 64546 265854
rect 64782 265618 64866 265854
rect 65102 265618 104546 265854
rect 104782 265618 104866 265854
rect 105102 265618 144546 265854
rect 144782 265618 144866 265854
rect 145102 265618 184546 265854
rect 184782 265618 184866 265854
rect 185102 265618 224546 265854
rect 224782 265618 224866 265854
rect 225102 265618 264546 265854
rect 264782 265618 264866 265854
rect 265102 265618 304546 265854
rect 304782 265618 304866 265854
rect 305102 265618 344546 265854
rect 344782 265618 344866 265854
rect 345102 265618 384546 265854
rect 384782 265618 384866 265854
rect 385102 265618 424546 265854
rect 424782 265618 424866 265854
rect 425102 265618 464546 265854
rect 464782 265618 464866 265854
rect 465102 265618 504546 265854
rect 504782 265618 504866 265854
rect 505102 265618 544546 265854
rect 544782 265618 544866 265854
rect 545102 265618 588222 265854
rect 588458 265618 588542 265854
rect 588778 265618 588810 265854
rect -4886 265586 588810 265618
rect -2966 262454 586890 262486
rect -2966 262218 -2934 262454
rect -2698 262218 -2614 262454
rect -2378 262218 20826 262454
rect 21062 262218 21146 262454
rect 21382 262218 60826 262454
rect 61062 262218 61146 262454
rect 61382 262218 100826 262454
rect 101062 262218 101146 262454
rect 101382 262218 140826 262454
rect 141382 262218 180826 262454
rect 181382 262218 220826 262454
rect 221382 262218 260826 262454
rect 261382 262218 300826 262454
rect 301382 262218 340826 262454
rect 341062 262218 341146 262454
rect 341382 262218 380826 262454
rect 381062 262218 381146 262454
rect 381382 262218 420826 262454
rect 421062 262218 421146 262454
rect 421382 262218 460826 262454
rect 461062 262218 461146 262454
rect 461382 262218 500826 262454
rect 501062 262218 501146 262454
rect 501382 262218 540826 262454
rect 541062 262218 541146 262454
rect 541382 262218 580826 262454
rect 581062 262218 581146 262454
rect 581382 262218 586302 262454
rect 586538 262218 586622 262454
rect 586858 262218 586890 262454
rect -2966 262134 586890 262218
rect -2966 261898 -2934 262134
rect -2698 261898 -2614 262134
rect -2378 261898 20826 262134
rect 21062 261898 21146 262134
rect 21382 261898 60826 262134
rect 61062 261898 61146 262134
rect 61382 261898 100826 262134
rect 101062 261898 101146 262134
rect 101382 261898 140826 262134
rect 141382 261898 180826 262134
rect 181382 261898 220826 262134
rect 221382 261898 260826 262134
rect 261382 261898 300826 262134
rect 301382 261898 340826 262134
rect 341062 261898 341146 262134
rect 341382 261898 380826 262134
rect 381062 261898 381146 262134
rect 381382 261898 420826 262134
rect 421062 261898 421146 262134
rect 421382 261898 460826 262134
rect 461062 261898 461146 262134
rect 461382 261898 500826 262134
rect 501062 261898 501146 262134
rect 501382 261898 540826 262134
rect 541062 261898 541146 262134
rect 541382 261898 580826 262134
rect 581062 261898 581146 262134
rect 581382 261898 586302 262134
rect 586538 261898 586622 262134
rect 586858 261898 586890 262134
rect -2966 261866 586890 261898
rect -8726 253614 592650 253646
rect -8726 253378 -7734 253614
rect -7498 253378 -7414 253614
rect -7178 253378 11986 253614
rect 12222 253378 12306 253614
rect 12542 253378 51986 253614
rect 52222 253378 52306 253614
rect 52542 253378 91986 253614
rect 92222 253378 92306 253614
rect 92542 253378 131986 253614
rect 132222 253378 132306 253614
rect 132542 253378 171986 253614
rect 172222 253378 172306 253614
rect 172542 253378 211986 253614
rect 212222 253378 212306 253614
rect 212542 253378 251986 253614
rect 252222 253378 252306 253614
rect 252542 253378 291986 253614
rect 292222 253378 292306 253614
rect 292542 253378 331986 253614
rect 332222 253378 332306 253614
rect 332542 253378 371986 253614
rect 372222 253378 372306 253614
rect 372542 253378 411986 253614
rect 412222 253378 412306 253614
rect 412542 253378 451986 253614
rect 452222 253378 452306 253614
rect 452542 253378 491986 253614
rect 492222 253378 492306 253614
rect 492542 253378 531986 253614
rect 532222 253378 532306 253614
rect 532542 253378 571986 253614
rect 572222 253378 572306 253614
rect 572542 253378 591102 253614
rect 591338 253378 591422 253614
rect 591658 253378 592650 253614
rect -8726 253294 592650 253378
rect -8726 253058 -7734 253294
rect -7498 253058 -7414 253294
rect -7178 253058 11986 253294
rect 12222 253058 12306 253294
rect 12542 253058 51986 253294
rect 52222 253058 52306 253294
rect 52542 253058 91986 253294
rect 92222 253058 92306 253294
rect 92542 253058 131986 253294
rect 132222 253058 132306 253294
rect 132542 253058 171986 253294
rect 172222 253058 172306 253294
rect 172542 253058 211986 253294
rect 212222 253058 212306 253294
rect 212542 253058 251986 253294
rect 252222 253058 252306 253294
rect 252542 253058 291986 253294
rect 292222 253058 292306 253294
rect 292542 253058 331986 253294
rect 332222 253058 332306 253294
rect 332542 253058 371986 253294
rect 372222 253058 372306 253294
rect 372542 253058 411986 253294
rect 412222 253058 412306 253294
rect 412542 253058 451986 253294
rect 452222 253058 452306 253294
rect 452542 253058 491986 253294
rect 492222 253058 492306 253294
rect 492542 253058 531986 253294
rect 532222 253058 532306 253294
rect 532542 253058 571986 253294
rect 572222 253058 572306 253294
rect 572542 253058 591102 253294
rect 591338 253058 591422 253294
rect 591658 253058 592650 253294
rect -8726 253026 592650 253058
rect -6806 249894 590730 249926
rect -6806 249658 -5814 249894
rect -5578 249658 -5494 249894
rect -5258 249658 8266 249894
rect 8502 249658 8586 249894
rect 8822 249658 48266 249894
rect 48502 249658 48586 249894
rect 48822 249658 88266 249894
rect 88502 249658 88586 249894
rect 88822 249658 128266 249894
rect 128502 249658 128586 249894
rect 128822 249658 168266 249894
rect 168502 249658 168586 249894
rect 168822 249658 208266 249894
rect 208502 249658 208586 249894
rect 208822 249658 248266 249894
rect 248502 249658 248586 249894
rect 248822 249658 288266 249894
rect 288502 249658 288586 249894
rect 288822 249658 328266 249894
rect 328502 249658 328586 249894
rect 328822 249658 368266 249894
rect 368502 249658 368586 249894
rect 368822 249658 408266 249894
rect 408502 249658 408586 249894
rect 408822 249658 448266 249894
rect 448502 249658 448586 249894
rect 448822 249658 488266 249894
rect 488502 249658 488586 249894
rect 488822 249658 528266 249894
rect 528502 249658 528586 249894
rect 528822 249658 568266 249894
rect 568502 249658 568586 249894
rect 568822 249658 589182 249894
rect 589418 249658 589502 249894
rect 589738 249658 590730 249894
rect -6806 249574 590730 249658
rect -6806 249338 -5814 249574
rect -5578 249338 -5494 249574
rect -5258 249338 8266 249574
rect 8502 249338 8586 249574
rect 8822 249338 48266 249574
rect 48502 249338 48586 249574
rect 48822 249338 88266 249574
rect 88502 249338 88586 249574
rect 88822 249338 128266 249574
rect 128502 249338 128586 249574
rect 128822 249338 168266 249574
rect 168502 249338 168586 249574
rect 168822 249338 208266 249574
rect 208502 249338 208586 249574
rect 208822 249338 248266 249574
rect 248502 249338 248586 249574
rect 248822 249338 288266 249574
rect 288502 249338 288586 249574
rect 288822 249338 328266 249574
rect 328502 249338 328586 249574
rect 328822 249338 368266 249574
rect 368502 249338 368586 249574
rect 368822 249338 408266 249574
rect 408502 249338 408586 249574
rect 408822 249338 448266 249574
rect 448502 249338 448586 249574
rect 448822 249338 488266 249574
rect 488502 249338 488586 249574
rect 488822 249338 528266 249574
rect 528502 249338 528586 249574
rect 528822 249338 568266 249574
rect 568502 249338 568586 249574
rect 568822 249338 589182 249574
rect 589418 249338 589502 249574
rect 589738 249338 590730 249574
rect -6806 249306 590730 249338
rect -4886 246174 588810 246206
rect -4886 245938 -3894 246174
rect -3658 245938 -3574 246174
rect -3338 245938 4546 246174
rect 4782 245938 4866 246174
rect 5102 245938 44546 246174
rect 44782 245938 44866 246174
rect 45102 245938 84546 246174
rect 84782 245938 84866 246174
rect 85102 245938 124546 246174
rect 124782 245938 124866 246174
rect 125102 245938 164546 246174
rect 164782 245938 164866 246174
rect 165102 245938 204546 246174
rect 204782 245938 204866 246174
rect 205102 245938 244546 246174
rect 244782 245938 244866 246174
rect 245102 245938 284546 246174
rect 284782 245938 284866 246174
rect 285102 245938 324546 246174
rect 324782 245938 324866 246174
rect 325102 245938 364546 246174
rect 364782 245938 364866 246174
rect 365102 245938 404546 246174
rect 404782 245938 404866 246174
rect 405102 245938 444546 246174
rect 444782 245938 444866 246174
rect 445102 245938 484546 246174
rect 484782 245938 484866 246174
rect 485102 245938 524546 246174
rect 524782 245938 524866 246174
rect 525102 245938 564546 246174
rect 564782 245938 564866 246174
rect 565102 245938 587262 246174
rect 587498 245938 587582 246174
rect 587818 245938 588810 246174
rect -4886 245854 588810 245938
rect -4886 245618 -3894 245854
rect -3658 245618 -3574 245854
rect -3338 245618 4546 245854
rect 4782 245618 4866 245854
rect 5102 245618 44546 245854
rect 44782 245618 44866 245854
rect 45102 245618 84546 245854
rect 84782 245618 84866 245854
rect 85102 245618 124546 245854
rect 124782 245618 124866 245854
rect 125102 245618 164546 245854
rect 164782 245618 164866 245854
rect 165102 245618 204546 245854
rect 204782 245618 204866 245854
rect 205102 245618 244546 245854
rect 244782 245618 244866 245854
rect 245102 245618 284546 245854
rect 284782 245618 284866 245854
rect 285102 245618 324546 245854
rect 324782 245618 324866 245854
rect 325102 245618 364546 245854
rect 364782 245618 364866 245854
rect 365102 245618 404546 245854
rect 404782 245618 404866 245854
rect 405102 245618 444546 245854
rect 444782 245618 444866 245854
rect 445102 245618 484546 245854
rect 484782 245618 484866 245854
rect 485102 245618 524546 245854
rect 524782 245618 524866 245854
rect 525102 245618 564546 245854
rect 564782 245618 564866 245854
rect 565102 245618 587262 245854
rect 587498 245618 587582 245854
rect 587818 245618 588810 245854
rect -4886 245586 588810 245618
rect -2966 242454 586890 242486
rect -2966 242218 -1974 242454
rect -1738 242218 -1654 242454
rect -1418 242218 826 242454
rect 1062 242218 1146 242454
rect 1382 242218 40826 242454
rect 41062 242218 41146 242454
rect 41382 242218 80826 242454
rect 81062 242218 81146 242454
rect 81382 242218 120826 242454
rect 121062 242218 121146 242454
rect 121382 242218 160826 242454
rect 161382 242218 200826 242454
rect 201382 242218 240826 242454
rect 241382 242218 280826 242454
rect 281382 242218 320826 242454
rect 321062 242218 321146 242454
rect 321382 242218 360826 242454
rect 361062 242218 361146 242454
rect 361382 242218 400826 242454
rect 401062 242218 401146 242454
rect 401382 242218 440826 242454
rect 441062 242218 441146 242454
rect 441382 242218 480826 242454
rect 481062 242218 481146 242454
rect 481382 242218 520826 242454
rect 521062 242218 521146 242454
rect 521382 242218 560826 242454
rect 561062 242218 561146 242454
rect 561382 242218 585342 242454
rect 585578 242218 585662 242454
rect 585898 242218 586890 242454
rect -2966 242134 586890 242218
rect -2966 241898 -1974 242134
rect -1738 241898 -1654 242134
rect -1418 241898 826 242134
rect 1062 241898 1146 242134
rect 1382 241898 40826 242134
rect 41062 241898 41146 242134
rect 41382 241898 80826 242134
rect 81062 241898 81146 242134
rect 81382 241898 120826 242134
rect 121062 241898 121146 242134
rect 121382 241898 160826 242134
rect 161382 241898 200826 242134
rect 201382 241898 240826 242134
rect 241382 241898 280826 242134
rect 281382 241898 320826 242134
rect 321062 241898 321146 242134
rect 321382 241898 360826 242134
rect 361062 241898 361146 242134
rect 361382 241898 400826 242134
rect 401062 241898 401146 242134
rect 401382 241898 440826 242134
rect 441062 241898 441146 242134
rect 441382 241898 480826 242134
rect 481062 241898 481146 242134
rect 481382 241898 520826 242134
rect 521062 241898 521146 242134
rect 521382 241898 560826 242134
rect 561062 241898 561146 242134
rect 561382 241898 585342 242134
rect 585578 241898 585662 242134
rect 585898 241898 586890 242134
rect -2966 241866 586890 241898
rect -8726 233614 592650 233646
rect -8726 233378 -8694 233614
rect -8458 233378 -8374 233614
rect -8138 233378 31986 233614
rect 32222 233378 32306 233614
rect 32542 233378 71986 233614
rect 72222 233378 72306 233614
rect 72542 233378 111986 233614
rect 112222 233378 112306 233614
rect 112542 233378 151986 233614
rect 152222 233378 152306 233614
rect 152542 233378 191986 233614
rect 192222 233378 192306 233614
rect 192542 233378 231986 233614
rect 232222 233378 232306 233614
rect 232542 233378 271986 233614
rect 272222 233378 272306 233614
rect 272542 233378 311986 233614
rect 312222 233378 312306 233614
rect 312542 233378 351986 233614
rect 352222 233378 352306 233614
rect 352542 233378 391986 233614
rect 392222 233378 392306 233614
rect 392542 233378 431986 233614
rect 432222 233378 432306 233614
rect 432542 233378 471986 233614
rect 472222 233378 472306 233614
rect 472542 233378 511986 233614
rect 512222 233378 512306 233614
rect 512542 233378 551986 233614
rect 552222 233378 552306 233614
rect 552542 233378 592062 233614
rect 592298 233378 592382 233614
rect 592618 233378 592650 233614
rect -8726 233294 592650 233378
rect -8726 233058 -8694 233294
rect -8458 233058 -8374 233294
rect -8138 233058 31986 233294
rect 32222 233058 32306 233294
rect 32542 233058 71986 233294
rect 72222 233058 72306 233294
rect 72542 233058 111986 233294
rect 112222 233058 112306 233294
rect 112542 233058 151986 233294
rect 152222 233058 152306 233294
rect 152542 233058 191986 233294
rect 192222 233058 192306 233294
rect 192542 233058 231986 233294
rect 232222 233058 232306 233294
rect 232542 233058 271986 233294
rect 272222 233058 272306 233294
rect 272542 233058 311986 233294
rect 312222 233058 312306 233294
rect 312542 233058 351986 233294
rect 352222 233058 352306 233294
rect 352542 233058 391986 233294
rect 392222 233058 392306 233294
rect 392542 233058 431986 233294
rect 432222 233058 432306 233294
rect 432542 233058 471986 233294
rect 472222 233058 472306 233294
rect 472542 233058 511986 233294
rect 512222 233058 512306 233294
rect 512542 233058 551986 233294
rect 552222 233058 552306 233294
rect 552542 233058 592062 233294
rect 592298 233058 592382 233294
rect 592618 233058 592650 233294
rect -8726 233026 592650 233058
rect -6806 229894 590730 229926
rect -6806 229658 -6774 229894
rect -6538 229658 -6454 229894
rect -6218 229658 28266 229894
rect 28502 229658 28586 229894
rect 28822 229658 68266 229894
rect 68502 229658 68586 229894
rect 68822 229658 108266 229894
rect 108502 229658 108586 229894
rect 108822 229658 148266 229894
rect 148502 229658 148586 229894
rect 148822 229658 188266 229894
rect 188502 229658 188586 229894
rect 188822 229658 228266 229894
rect 228502 229658 228586 229894
rect 228822 229658 268266 229894
rect 268502 229658 268586 229894
rect 268822 229658 308266 229894
rect 308502 229658 308586 229894
rect 308822 229658 348266 229894
rect 348502 229658 348586 229894
rect 348822 229658 388266 229894
rect 388502 229658 388586 229894
rect 388822 229658 428266 229894
rect 428502 229658 428586 229894
rect 428822 229658 468266 229894
rect 468502 229658 468586 229894
rect 468822 229658 508266 229894
rect 508502 229658 508586 229894
rect 508822 229658 548266 229894
rect 548502 229658 548586 229894
rect 548822 229658 590142 229894
rect 590378 229658 590462 229894
rect 590698 229658 590730 229894
rect -6806 229574 590730 229658
rect -6806 229338 -6774 229574
rect -6538 229338 -6454 229574
rect -6218 229338 28266 229574
rect 28502 229338 28586 229574
rect 28822 229338 68266 229574
rect 68502 229338 68586 229574
rect 68822 229338 108266 229574
rect 108502 229338 108586 229574
rect 108822 229338 148266 229574
rect 148502 229338 148586 229574
rect 148822 229338 188266 229574
rect 188502 229338 188586 229574
rect 188822 229338 228266 229574
rect 228502 229338 228586 229574
rect 228822 229338 268266 229574
rect 268502 229338 268586 229574
rect 268822 229338 308266 229574
rect 308502 229338 308586 229574
rect 308822 229338 348266 229574
rect 348502 229338 348586 229574
rect 348822 229338 388266 229574
rect 388502 229338 388586 229574
rect 388822 229338 428266 229574
rect 428502 229338 428586 229574
rect 428822 229338 468266 229574
rect 468502 229338 468586 229574
rect 468822 229338 508266 229574
rect 508502 229338 508586 229574
rect 508822 229338 548266 229574
rect 548502 229338 548586 229574
rect 548822 229338 590142 229574
rect 590378 229338 590462 229574
rect 590698 229338 590730 229574
rect -6806 229306 590730 229338
rect -4886 226174 588810 226206
rect -4886 225938 -4854 226174
rect -4618 225938 -4534 226174
rect -4298 225938 24546 226174
rect 24782 225938 24866 226174
rect 25102 225938 64546 226174
rect 64782 225938 64866 226174
rect 65102 225938 104546 226174
rect 104782 225938 104866 226174
rect 105102 225938 144546 226174
rect 144782 225938 144866 226174
rect 145102 225938 184546 226174
rect 184782 225938 184866 226174
rect 185102 225938 224546 226174
rect 224782 225938 224866 226174
rect 225102 225938 264546 226174
rect 264782 225938 264866 226174
rect 265102 225938 304546 226174
rect 304782 225938 304866 226174
rect 305102 225938 344546 226174
rect 344782 225938 344866 226174
rect 345102 225938 384546 226174
rect 384782 225938 384866 226174
rect 385102 225938 424546 226174
rect 424782 225938 424866 226174
rect 425102 225938 464546 226174
rect 464782 225938 464866 226174
rect 465102 225938 504546 226174
rect 504782 225938 504866 226174
rect 505102 225938 544546 226174
rect 544782 225938 544866 226174
rect 545102 225938 588222 226174
rect 588458 225938 588542 226174
rect 588778 225938 588810 226174
rect -4886 225854 588810 225938
rect -4886 225618 -4854 225854
rect -4618 225618 -4534 225854
rect -4298 225618 24546 225854
rect 24782 225618 24866 225854
rect 25102 225618 64546 225854
rect 64782 225618 64866 225854
rect 65102 225618 104546 225854
rect 104782 225618 104866 225854
rect 105102 225618 144546 225854
rect 144782 225618 144866 225854
rect 145102 225618 184546 225854
rect 184782 225618 184866 225854
rect 185102 225618 224546 225854
rect 224782 225618 224866 225854
rect 225102 225618 264546 225854
rect 264782 225618 264866 225854
rect 265102 225618 304546 225854
rect 304782 225618 304866 225854
rect 305102 225618 344546 225854
rect 344782 225618 344866 225854
rect 345102 225618 384546 225854
rect 384782 225618 384866 225854
rect 385102 225618 424546 225854
rect 424782 225618 424866 225854
rect 425102 225618 464546 225854
rect 464782 225618 464866 225854
rect 465102 225618 504546 225854
rect 504782 225618 504866 225854
rect 505102 225618 544546 225854
rect 544782 225618 544866 225854
rect 545102 225618 588222 225854
rect 588458 225618 588542 225854
rect 588778 225618 588810 225854
rect -4886 225586 588810 225618
rect -2966 222454 586890 222486
rect -2966 222218 -2934 222454
rect -2698 222218 -2614 222454
rect -2378 222218 20826 222454
rect 21062 222218 21146 222454
rect 21382 222218 60826 222454
rect 61062 222218 61146 222454
rect 61382 222218 100826 222454
rect 101062 222218 101146 222454
rect 101382 222218 140826 222454
rect 141382 222218 180826 222454
rect 181382 222218 220826 222454
rect 221382 222218 260826 222454
rect 261382 222218 300826 222454
rect 301382 222218 340826 222454
rect 341062 222218 341146 222454
rect 341382 222218 380826 222454
rect 381062 222218 381146 222454
rect 381382 222218 420826 222454
rect 421062 222218 421146 222454
rect 421382 222218 460826 222454
rect 461062 222218 461146 222454
rect 461382 222218 500826 222454
rect 501062 222218 501146 222454
rect 501382 222218 540826 222454
rect 541062 222218 541146 222454
rect 541382 222218 580826 222454
rect 581062 222218 581146 222454
rect 581382 222218 586302 222454
rect 586538 222218 586622 222454
rect 586858 222218 586890 222454
rect -2966 222134 586890 222218
rect -2966 221898 -2934 222134
rect -2698 221898 -2614 222134
rect -2378 221898 20826 222134
rect 21062 221898 21146 222134
rect 21382 221898 60826 222134
rect 61062 221898 61146 222134
rect 61382 221898 100826 222134
rect 101062 221898 101146 222134
rect 101382 221898 140826 222134
rect 141382 221898 180826 222134
rect 181382 221898 220826 222134
rect 221382 221898 260826 222134
rect 261382 221898 300826 222134
rect 301382 221898 340826 222134
rect 341062 221898 341146 222134
rect 341382 221898 380826 222134
rect 381062 221898 381146 222134
rect 381382 221898 420826 222134
rect 421062 221898 421146 222134
rect 421382 221898 460826 222134
rect 461062 221898 461146 222134
rect 461382 221898 500826 222134
rect 501062 221898 501146 222134
rect 501382 221898 540826 222134
rect 541062 221898 541146 222134
rect 541382 221898 580826 222134
rect 581062 221898 581146 222134
rect 581382 221898 586302 222134
rect 586538 221898 586622 222134
rect 586858 221898 586890 222134
rect -2966 221866 586890 221898
rect -8726 213614 592650 213646
rect -8726 213378 -7734 213614
rect -7498 213378 -7414 213614
rect -7178 213378 11986 213614
rect 12222 213378 12306 213614
rect 12542 213378 51986 213614
rect 52222 213378 52306 213614
rect 52542 213378 91986 213614
rect 92222 213378 92306 213614
rect 92542 213378 131986 213614
rect 132222 213378 132306 213614
rect 132542 213378 171986 213614
rect 172222 213378 172306 213614
rect 172542 213378 211986 213614
rect 212222 213378 212306 213614
rect 212542 213378 251986 213614
rect 252222 213378 252306 213614
rect 252542 213378 291986 213614
rect 292222 213378 292306 213614
rect 292542 213378 331986 213614
rect 332222 213378 332306 213614
rect 332542 213378 371986 213614
rect 372222 213378 372306 213614
rect 372542 213378 411986 213614
rect 412222 213378 412306 213614
rect 412542 213378 451986 213614
rect 452222 213378 452306 213614
rect 452542 213378 491986 213614
rect 492222 213378 492306 213614
rect 492542 213378 531986 213614
rect 532222 213378 532306 213614
rect 532542 213378 571986 213614
rect 572222 213378 572306 213614
rect 572542 213378 591102 213614
rect 591338 213378 591422 213614
rect 591658 213378 592650 213614
rect -8726 213294 592650 213378
rect -8726 213058 -7734 213294
rect -7498 213058 -7414 213294
rect -7178 213058 11986 213294
rect 12222 213058 12306 213294
rect 12542 213058 51986 213294
rect 52222 213058 52306 213294
rect 52542 213058 91986 213294
rect 92222 213058 92306 213294
rect 92542 213058 131986 213294
rect 132222 213058 132306 213294
rect 132542 213058 171986 213294
rect 172222 213058 172306 213294
rect 172542 213058 211986 213294
rect 212222 213058 212306 213294
rect 212542 213058 251986 213294
rect 252222 213058 252306 213294
rect 252542 213058 291986 213294
rect 292222 213058 292306 213294
rect 292542 213058 331986 213294
rect 332222 213058 332306 213294
rect 332542 213058 371986 213294
rect 372222 213058 372306 213294
rect 372542 213058 411986 213294
rect 412222 213058 412306 213294
rect 412542 213058 451986 213294
rect 452222 213058 452306 213294
rect 452542 213058 491986 213294
rect 492222 213058 492306 213294
rect 492542 213058 531986 213294
rect 532222 213058 532306 213294
rect 532542 213058 571986 213294
rect 572222 213058 572306 213294
rect 572542 213058 591102 213294
rect 591338 213058 591422 213294
rect 591658 213058 592650 213294
rect -8726 213026 592650 213058
rect -6806 209894 590730 209926
rect -6806 209658 -5814 209894
rect -5578 209658 -5494 209894
rect -5258 209658 8266 209894
rect 8502 209658 8586 209894
rect 8822 209658 48266 209894
rect 48502 209658 48586 209894
rect 48822 209658 88266 209894
rect 88502 209658 88586 209894
rect 88822 209658 128266 209894
rect 128502 209658 128586 209894
rect 128822 209658 168266 209894
rect 168502 209658 168586 209894
rect 168822 209658 208266 209894
rect 208502 209658 208586 209894
rect 208822 209658 248266 209894
rect 248502 209658 248586 209894
rect 248822 209658 288266 209894
rect 288502 209658 288586 209894
rect 288822 209658 328266 209894
rect 328502 209658 328586 209894
rect 328822 209658 368266 209894
rect 368502 209658 368586 209894
rect 368822 209658 408266 209894
rect 408502 209658 408586 209894
rect 408822 209658 448266 209894
rect 448502 209658 448586 209894
rect 448822 209658 488266 209894
rect 488502 209658 488586 209894
rect 488822 209658 528266 209894
rect 528502 209658 528586 209894
rect 528822 209658 568266 209894
rect 568502 209658 568586 209894
rect 568822 209658 589182 209894
rect 589418 209658 589502 209894
rect 589738 209658 590730 209894
rect -6806 209574 590730 209658
rect -6806 209338 -5814 209574
rect -5578 209338 -5494 209574
rect -5258 209338 8266 209574
rect 8502 209338 8586 209574
rect 8822 209338 48266 209574
rect 48502 209338 48586 209574
rect 48822 209338 88266 209574
rect 88502 209338 88586 209574
rect 88822 209338 128266 209574
rect 128502 209338 128586 209574
rect 128822 209338 168266 209574
rect 168502 209338 168586 209574
rect 168822 209338 208266 209574
rect 208502 209338 208586 209574
rect 208822 209338 248266 209574
rect 248502 209338 248586 209574
rect 248822 209338 288266 209574
rect 288502 209338 288586 209574
rect 288822 209338 328266 209574
rect 328502 209338 328586 209574
rect 328822 209338 368266 209574
rect 368502 209338 368586 209574
rect 368822 209338 408266 209574
rect 408502 209338 408586 209574
rect 408822 209338 448266 209574
rect 448502 209338 448586 209574
rect 448822 209338 488266 209574
rect 488502 209338 488586 209574
rect 488822 209338 528266 209574
rect 528502 209338 528586 209574
rect 528822 209338 568266 209574
rect 568502 209338 568586 209574
rect 568822 209338 589182 209574
rect 589418 209338 589502 209574
rect 589738 209338 590730 209574
rect -6806 209306 590730 209338
rect -4886 206174 588810 206206
rect -4886 205938 -3894 206174
rect -3658 205938 -3574 206174
rect -3338 205938 4546 206174
rect 4782 205938 4866 206174
rect 5102 205938 44546 206174
rect 44782 205938 44866 206174
rect 45102 205938 84546 206174
rect 84782 205938 84866 206174
rect 85102 205938 124546 206174
rect 124782 205938 124866 206174
rect 125102 205938 164546 206174
rect 164782 205938 164866 206174
rect 165102 205938 204546 206174
rect 204782 205938 204866 206174
rect 205102 205938 244546 206174
rect 244782 205938 244866 206174
rect 245102 205938 284546 206174
rect 284782 205938 284866 206174
rect 285102 205938 324546 206174
rect 324782 205938 324866 206174
rect 325102 205938 364546 206174
rect 364782 205938 364866 206174
rect 365102 205938 404546 206174
rect 404782 205938 404866 206174
rect 405102 205938 444546 206174
rect 444782 205938 444866 206174
rect 445102 205938 484546 206174
rect 484782 205938 484866 206174
rect 485102 205938 524546 206174
rect 524782 205938 524866 206174
rect 525102 205938 564546 206174
rect 564782 205938 564866 206174
rect 565102 205938 587262 206174
rect 587498 205938 587582 206174
rect 587818 205938 588810 206174
rect -4886 205854 588810 205938
rect -4886 205618 -3894 205854
rect -3658 205618 -3574 205854
rect -3338 205618 4546 205854
rect 4782 205618 4866 205854
rect 5102 205618 44546 205854
rect 44782 205618 44866 205854
rect 45102 205618 84546 205854
rect 84782 205618 84866 205854
rect 85102 205618 124546 205854
rect 124782 205618 124866 205854
rect 125102 205618 164546 205854
rect 164782 205618 164866 205854
rect 165102 205618 204546 205854
rect 204782 205618 204866 205854
rect 205102 205618 244546 205854
rect 244782 205618 244866 205854
rect 245102 205618 284546 205854
rect 284782 205618 284866 205854
rect 285102 205618 324546 205854
rect 324782 205618 324866 205854
rect 325102 205618 364546 205854
rect 364782 205618 364866 205854
rect 365102 205618 404546 205854
rect 404782 205618 404866 205854
rect 405102 205618 444546 205854
rect 444782 205618 444866 205854
rect 445102 205618 484546 205854
rect 484782 205618 484866 205854
rect 485102 205618 524546 205854
rect 524782 205618 524866 205854
rect 525102 205618 564546 205854
rect 564782 205618 564866 205854
rect 565102 205618 587262 205854
rect 587498 205618 587582 205854
rect 587818 205618 588810 205854
rect -4886 205586 588810 205618
rect -2966 202454 586890 202486
rect -2966 202218 -1974 202454
rect -1738 202218 -1654 202454
rect -1418 202218 826 202454
rect 1062 202218 1146 202454
rect 1382 202218 40826 202454
rect 41062 202218 41146 202454
rect 41382 202218 80826 202454
rect 81062 202218 81146 202454
rect 81382 202218 120826 202454
rect 121062 202218 121146 202454
rect 121382 202218 160826 202454
rect 161382 202218 200826 202454
rect 201382 202218 240826 202454
rect 241382 202218 280826 202454
rect 281382 202218 320826 202454
rect 321062 202218 321146 202454
rect 321382 202218 360826 202454
rect 361062 202218 361146 202454
rect 361382 202218 400826 202454
rect 401062 202218 401146 202454
rect 401382 202218 440826 202454
rect 441062 202218 441146 202454
rect 441382 202218 480826 202454
rect 481062 202218 481146 202454
rect 481382 202218 520826 202454
rect 521062 202218 521146 202454
rect 521382 202218 560826 202454
rect 561062 202218 561146 202454
rect 561382 202218 585342 202454
rect 585578 202218 585662 202454
rect 585898 202218 586890 202454
rect -2966 202134 586890 202218
rect -2966 201898 -1974 202134
rect -1738 201898 -1654 202134
rect -1418 201898 826 202134
rect 1062 201898 1146 202134
rect 1382 201898 40826 202134
rect 41062 201898 41146 202134
rect 41382 201898 80826 202134
rect 81062 201898 81146 202134
rect 81382 201898 120826 202134
rect 121062 201898 121146 202134
rect 121382 201898 160826 202134
rect 161382 201898 200826 202134
rect 201382 201898 240826 202134
rect 241382 201898 280826 202134
rect 281382 201898 320826 202134
rect 321062 201898 321146 202134
rect 321382 201898 360826 202134
rect 361062 201898 361146 202134
rect 361382 201898 400826 202134
rect 401062 201898 401146 202134
rect 401382 201898 440826 202134
rect 441062 201898 441146 202134
rect 441382 201898 480826 202134
rect 481062 201898 481146 202134
rect 481382 201898 520826 202134
rect 521062 201898 521146 202134
rect 521382 201898 560826 202134
rect 561062 201898 561146 202134
rect 561382 201898 585342 202134
rect 585578 201898 585662 202134
rect 585898 201898 586890 202134
rect -2966 201866 586890 201898
rect -8726 193614 592650 193646
rect -8726 193378 -8694 193614
rect -8458 193378 -8374 193614
rect -8138 193378 31986 193614
rect 32222 193378 32306 193614
rect 32542 193378 71986 193614
rect 72222 193378 72306 193614
rect 72542 193378 111986 193614
rect 112222 193378 112306 193614
rect 112542 193378 151986 193614
rect 152222 193378 152306 193614
rect 152542 193378 191986 193614
rect 192222 193378 192306 193614
rect 192542 193378 231986 193614
rect 232222 193378 232306 193614
rect 232542 193378 271986 193614
rect 272222 193378 272306 193614
rect 272542 193378 311986 193614
rect 312222 193378 312306 193614
rect 312542 193378 351986 193614
rect 352222 193378 352306 193614
rect 352542 193378 391986 193614
rect 392222 193378 392306 193614
rect 392542 193378 431986 193614
rect 432222 193378 432306 193614
rect 432542 193378 471986 193614
rect 472222 193378 472306 193614
rect 472542 193378 511986 193614
rect 512222 193378 512306 193614
rect 512542 193378 551986 193614
rect 552222 193378 552306 193614
rect 552542 193378 592062 193614
rect 592298 193378 592382 193614
rect 592618 193378 592650 193614
rect -8726 193294 592650 193378
rect -8726 193058 -8694 193294
rect -8458 193058 -8374 193294
rect -8138 193058 31986 193294
rect 32222 193058 32306 193294
rect 32542 193058 71986 193294
rect 72222 193058 72306 193294
rect 72542 193058 111986 193294
rect 112222 193058 112306 193294
rect 112542 193058 151986 193294
rect 152222 193058 152306 193294
rect 152542 193058 191986 193294
rect 192222 193058 192306 193294
rect 192542 193058 231986 193294
rect 232222 193058 232306 193294
rect 232542 193058 271986 193294
rect 272222 193058 272306 193294
rect 272542 193058 311986 193294
rect 312222 193058 312306 193294
rect 312542 193058 351986 193294
rect 352222 193058 352306 193294
rect 352542 193058 391986 193294
rect 392222 193058 392306 193294
rect 392542 193058 431986 193294
rect 432222 193058 432306 193294
rect 432542 193058 471986 193294
rect 472222 193058 472306 193294
rect 472542 193058 511986 193294
rect 512222 193058 512306 193294
rect 512542 193058 551986 193294
rect 552222 193058 552306 193294
rect 552542 193058 592062 193294
rect 592298 193058 592382 193294
rect 592618 193058 592650 193294
rect -8726 193026 592650 193058
rect -6806 189894 590730 189926
rect -6806 189658 -6774 189894
rect -6538 189658 -6454 189894
rect -6218 189658 28266 189894
rect 28502 189658 28586 189894
rect 28822 189658 68266 189894
rect 68502 189658 68586 189894
rect 68822 189658 108266 189894
rect 108502 189658 108586 189894
rect 108822 189658 148266 189894
rect 148502 189658 148586 189894
rect 148822 189658 188266 189894
rect 188502 189658 188586 189894
rect 188822 189658 228266 189894
rect 228502 189658 228586 189894
rect 228822 189658 268266 189894
rect 268502 189658 268586 189894
rect 268822 189658 308266 189894
rect 308502 189658 308586 189894
rect 308822 189658 348266 189894
rect 348502 189658 348586 189894
rect 348822 189658 388266 189894
rect 388502 189658 388586 189894
rect 388822 189658 428266 189894
rect 428502 189658 428586 189894
rect 428822 189658 468266 189894
rect 468502 189658 468586 189894
rect 468822 189658 508266 189894
rect 508502 189658 508586 189894
rect 508822 189658 548266 189894
rect 548502 189658 548586 189894
rect 548822 189658 590142 189894
rect 590378 189658 590462 189894
rect 590698 189658 590730 189894
rect -6806 189574 590730 189658
rect -6806 189338 -6774 189574
rect -6538 189338 -6454 189574
rect -6218 189338 28266 189574
rect 28502 189338 28586 189574
rect 28822 189338 68266 189574
rect 68502 189338 68586 189574
rect 68822 189338 108266 189574
rect 108502 189338 108586 189574
rect 108822 189338 148266 189574
rect 148502 189338 148586 189574
rect 148822 189338 188266 189574
rect 188502 189338 188586 189574
rect 188822 189338 228266 189574
rect 228502 189338 228586 189574
rect 228822 189338 268266 189574
rect 268502 189338 268586 189574
rect 268822 189338 308266 189574
rect 308502 189338 308586 189574
rect 308822 189338 348266 189574
rect 348502 189338 348586 189574
rect 348822 189338 388266 189574
rect 388502 189338 388586 189574
rect 388822 189338 428266 189574
rect 428502 189338 428586 189574
rect 428822 189338 468266 189574
rect 468502 189338 468586 189574
rect 468822 189338 508266 189574
rect 508502 189338 508586 189574
rect 508822 189338 548266 189574
rect 548502 189338 548586 189574
rect 548822 189338 590142 189574
rect 590378 189338 590462 189574
rect 590698 189338 590730 189574
rect -6806 189306 590730 189338
rect -4886 186174 588810 186206
rect -4886 185938 -4854 186174
rect -4618 185938 -4534 186174
rect -4298 185938 24546 186174
rect 24782 185938 24866 186174
rect 25102 185938 64546 186174
rect 64782 185938 64866 186174
rect 65102 185938 104546 186174
rect 104782 185938 104866 186174
rect 105102 185938 144546 186174
rect 144782 185938 144866 186174
rect 145102 185938 184546 186174
rect 184782 185938 184866 186174
rect 185102 185938 224546 186174
rect 224782 185938 224866 186174
rect 225102 185938 264546 186174
rect 264782 185938 264866 186174
rect 265102 185938 304546 186174
rect 304782 185938 304866 186174
rect 305102 185938 344546 186174
rect 344782 185938 344866 186174
rect 345102 185938 384546 186174
rect 384782 185938 384866 186174
rect 385102 185938 424546 186174
rect 424782 185938 424866 186174
rect 425102 185938 464546 186174
rect 464782 185938 464866 186174
rect 465102 185938 504546 186174
rect 504782 185938 504866 186174
rect 505102 185938 544546 186174
rect 544782 185938 544866 186174
rect 545102 185938 588222 186174
rect 588458 185938 588542 186174
rect 588778 185938 588810 186174
rect -4886 185854 588810 185938
rect -4886 185618 -4854 185854
rect -4618 185618 -4534 185854
rect -4298 185618 24546 185854
rect 24782 185618 24866 185854
rect 25102 185618 64546 185854
rect 64782 185618 64866 185854
rect 65102 185618 104546 185854
rect 104782 185618 104866 185854
rect 105102 185618 144546 185854
rect 144782 185618 144866 185854
rect 145102 185618 184546 185854
rect 184782 185618 184866 185854
rect 185102 185618 224546 185854
rect 224782 185618 224866 185854
rect 225102 185618 264546 185854
rect 264782 185618 264866 185854
rect 265102 185618 304546 185854
rect 304782 185618 304866 185854
rect 305102 185618 344546 185854
rect 344782 185618 344866 185854
rect 345102 185618 384546 185854
rect 384782 185618 384866 185854
rect 385102 185618 424546 185854
rect 424782 185618 424866 185854
rect 425102 185618 464546 185854
rect 464782 185618 464866 185854
rect 465102 185618 504546 185854
rect 504782 185618 504866 185854
rect 505102 185618 544546 185854
rect 544782 185618 544866 185854
rect 545102 185618 588222 185854
rect 588458 185618 588542 185854
rect 588778 185618 588810 185854
rect -4886 185586 588810 185618
rect -2966 182454 586890 182486
rect -2966 182218 -2934 182454
rect -2698 182218 -2614 182454
rect -2378 182218 20826 182454
rect 21062 182218 21146 182454
rect 21382 182218 60826 182454
rect 61062 182218 61146 182454
rect 61382 182218 100826 182454
rect 101062 182218 101146 182454
rect 101382 182218 140826 182454
rect 141382 182218 180826 182454
rect 181382 182218 220826 182454
rect 221382 182218 260826 182454
rect 261382 182218 300826 182454
rect 301382 182218 340826 182454
rect 341062 182218 341146 182454
rect 341382 182218 380826 182454
rect 381062 182218 381146 182454
rect 381382 182218 420826 182454
rect 421062 182218 421146 182454
rect 421382 182218 460826 182454
rect 461062 182218 461146 182454
rect 461382 182218 500826 182454
rect 501062 182218 501146 182454
rect 501382 182218 540826 182454
rect 541062 182218 541146 182454
rect 541382 182218 580826 182454
rect 581062 182218 581146 182454
rect 581382 182218 586302 182454
rect 586538 182218 586622 182454
rect 586858 182218 586890 182454
rect -2966 182134 586890 182218
rect -2966 181898 -2934 182134
rect -2698 181898 -2614 182134
rect -2378 181898 20826 182134
rect 21062 181898 21146 182134
rect 21382 181898 60826 182134
rect 61062 181898 61146 182134
rect 61382 181898 100826 182134
rect 101062 181898 101146 182134
rect 101382 181898 140826 182134
rect 141382 181898 180826 182134
rect 181382 181898 220826 182134
rect 221382 181898 260826 182134
rect 261382 181898 300826 182134
rect 301382 181898 340826 182134
rect 341062 181898 341146 182134
rect 341382 181898 380826 182134
rect 381062 181898 381146 182134
rect 381382 181898 420826 182134
rect 421062 181898 421146 182134
rect 421382 181898 460826 182134
rect 461062 181898 461146 182134
rect 461382 181898 500826 182134
rect 501062 181898 501146 182134
rect 501382 181898 540826 182134
rect 541062 181898 541146 182134
rect 541382 181898 580826 182134
rect 581062 181898 581146 182134
rect 581382 181898 586302 182134
rect 586538 181898 586622 182134
rect 586858 181898 586890 182134
rect -2966 181866 586890 181898
rect -8726 173614 592650 173646
rect -8726 173378 -7734 173614
rect -7498 173378 -7414 173614
rect -7178 173378 11986 173614
rect 12222 173378 12306 173614
rect 12542 173378 51986 173614
rect 52222 173378 52306 173614
rect 52542 173378 91986 173614
rect 92222 173378 92306 173614
rect 92542 173378 131986 173614
rect 132222 173378 132306 173614
rect 132542 173378 171986 173614
rect 172222 173378 172306 173614
rect 172542 173378 211986 173614
rect 212222 173378 212306 173614
rect 212542 173378 251986 173614
rect 252222 173378 252306 173614
rect 252542 173378 291986 173614
rect 292222 173378 292306 173614
rect 292542 173378 331986 173614
rect 332222 173378 332306 173614
rect 332542 173378 371986 173614
rect 372222 173378 372306 173614
rect 372542 173378 411986 173614
rect 412222 173378 412306 173614
rect 412542 173378 451986 173614
rect 452222 173378 452306 173614
rect 452542 173378 491986 173614
rect 492222 173378 492306 173614
rect 492542 173378 531986 173614
rect 532222 173378 532306 173614
rect 532542 173378 571986 173614
rect 572222 173378 572306 173614
rect 572542 173378 591102 173614
rect 591338 173378 591422 173614
rect 591658 173378 592650 173614
rect -8726 173294 592650 173378
rect -8726 173058 -7734 173294
rect -7498 173058 -7414 173294
rect -7178 173058 11986 173294
rect 12222 173058 12306 173294
rect 12542 173058 51986 173294
rect 52222 173058 52306 173294
rect 52542 173058 91986 173294
rect 92222 173058 92306 173294
rect 92542 173058 131986 173294
rect 132222 173058 132306 173294
rect 132542 173058 171986 173294
rect 172222 173058 172306 173294
rect 172542 173058 211986 173294
rect 212222 173058 212306 173294
rect 212542 173058 251986 173294
rect 252222 173058 252306 173294
rect 252542 173058 291986 173294
rect 292222 173058 292306 173294
rect 292542 173058 331986 173294
rect 332222 173058 332306 173294
rect 332542 173058 371986 173294
rect 372222 173058 372306 173294
rect 372542 173058 411986 173294
rect 412222 173058 412306 173294
rect 412542 173058 451986 173294
rect 452222 173058 452306 173294
rect 452542 173058 491986 173294
rect 492222 173058 492306 173294
rect 492542 173058 531986 173294
rect 532222 173058 532306 173294
rect 532542 173058 571986 173294
rect 572222 173058 572306 173294
rect 572542 173058 591102 173294
rect 591338 173058 591422 173294
rect 591658 173058 592650 173294
rect -8726 173026 592650 173058
rect -6806 169894 590730 169926
rect -6806 169658 -5814 169894
rect -5578 169658 -5494 169894
rect -5258 169658 8266 169894
rect 8502 169658 8586 169894
rect 8822 169658 48266 169894
rect 48502 169658 48586 169894
rect 48822 169658 88266 169894
rect 88502 169658 88586 169894
rect 88822 169658 128266 169894
rect 128502 169658 128586 169894
rect 128822 169658 168266 169894
rect 168502 169658 168586 169894
rect 168822 169658 208266 169894
rect 208502 169658 208586 169894
rect 208822 169658 248266 169894
rect 248502 169658 248586 169894
rect 248822 169658 288266 169894
rect 288502 169658 288586 169894
rect 288822 169658 328266 169894
rect 328502 169658 328586 169894
rect 328822 169658 368266 169894
rect 368502 169658 368586 169894
rect 368822 169658 408266 169894
rect 408502 169658 408586 169894
rect 408822 169658 448266 169894
rect 448502 169658 448586 169894
rect 448822 169658 488266 169894
rect 488502 169658 488586 169894
rect 488822 169658 528266 169894
rect 528502 169658 528586 169894
rect 528822 169658 568266 169894
rect 568502 169658 568586 169894
rect 568822 169658 589182 169894
rect 589418 169658 589502 169894
rect 589738 169658 590730 169894
rect -6806 169574 590730 169658
rect -6806 169338 -5814 169574
rect -5578 169338 -5494 169574
rect -5258 169338 8266 169574
rect 8502 169338 8586 169574
rect 8822 169338 48266 169574
rect 48502 169338 48586 169574
rect 48822 169338 88266 169574
rect 88502 169338 88586 169574
rect 88822 169338 128266 169574
rect 128502 169338 128586 169574
rect 128822 169338 168266 169574
rect 168502 169338 168586 169574
rect 168822 169338 208266 169574
rect 208502 169338 208586 169574
rect 208822 169338 248266 169574
rect 248502 169338 248586 169574
rect 248822 169338 288266 169574
rect 288502 169338 288586 169574
rect 288822 169338 328266 169574
rect 328502 169338 328586 169574
rect 328822 169338 368266 169574
rect 368502 169338 368586 169574
rect 368822 169338 408266 169574
rect 408502 169338 408586 169574
rect 408822 169338 448266 169574
rect 448502 169338 448586 169574
rect 448822 169338 488266 169574
rect 488502 169338 488586 169574
rect 488822 169338 528266 169574
rect 528502 169338 528586 169574
rect 528822 169338 568266 169574
rect 568502 169338 568586 169574
rect 568822 169338 589182 169574
rect 589418 169338 589502 169574
rect 589738 169338 590730 169574
rect -6806 169306 590730 169338
rect -4886 166174 588810 166206
rect -4886 165938 -3894 166174
rect -3658 165938 -3574 166174
rect -3338 165938 4546 166174
rect 4782 165938 4866 166174
rect 5102 165938 44546 166174
rect 44782 165938 44866 166174
rect 45102 165938 84546 166174
rect 84782 165938 84866 166174
rect 85102 165938 124546 166174
rect 124782 165938 124866 166174
rect 125102 165938 164546 166174
rect 164782 165938 164866 166174
rect 165102 165938 204546 166174
rect 204782 165938 204866 166174
rect 205102 165938 244546 166174
rect 244782 165938 244866 166174
rect 245102 165938 284546 166174
rect 284782 165938 284866 166174
rect 285102 165938 324546 166174
rect 324782 165938 324866 166174
rect 325102 165938 364546 166174
rect 364782 165938 364866 166174
rect 365102 165938 404546 166174
rect 404782 165938 404866 166174
rect 405102 165938 444546 166174
rect 444782 165938 444866 166174
rect 445102 165938 484546 166174
rect 484782 165938 484866 166174
rect 485102 165938 524546 166174
rect 524782 165938 524866 166174
rect 525102 165938 564546 166174
rect 564782 165938 564866 166174
rect 565102 165938 587262 166174
rect 587498 165938 587582 166174
rect 587818 165938 588810 166174
rect -4886 165854 588810 165938
rect -4886 165618 -3894 165854
rect -3658 165618 -3574 165854
rect -3338 165618 4546 165854
rect 4782 165618 4866 165854
rect 5102 165618 44546 165854
rect 44782 165618 44866 165854
rect 45102 165618 84546 165854
rect 84782 165618 84866 165854
rect 85102 165618 124546 165854
rect 124782 165618 124866 165854
rect 125102 165618 164546 165854
rect 164782 165618 164866 165854
rect 165102 165618 204546 165854
rect 204782 165618 204866 165854
rect 205102 165618 244546 165854
rect 244782 165618 244866 165854
rect 245102 165618 284546 165854
rect 284782 165618 284866 165854
rect 285102 165618 324546 165854
rect 324782 165618 324866 165854
rect 325102 165618 364546 165854
rect 364782 165618 364866 165854
rect 365102 165618 404546 165854
rect 404782 165618 404866 165854
rect 405102 165618 444546 165854
rect 444782 165618 444866 165854
rect 445102 165618 484546 165854
rect 484782 165618 484866 165854
rect 485102 165618 524546 165854
rect 524782 165618 524866 165854
rect 525102 165618 564546 165854
rect 564782 165618 564866 165854
rect 565102 165618 587262 165854
rect 587498 165618 587582 165854
rect 587818 165618 588810 165854
rect -4886 165586 588810 165618
rect -2966 162454 586890 162486
rect -2966 162218 -1974 162454
rect -1738 162218 -1654 162454
rect -1418 162218 826 162454
rect 1062 162218 1146 162454
rect 1382 162218 40826 162454
rect 41062 162218 41146 162454
rect 41382 162218 80826 162454
rect 81062 162218 81146 162454
rect 81382 162218 120826 162454
rect 121062 162218 121146 162454
rect 121382 162218 160826 162454
rect 161382 162218 200826 162454
rect 201382 162218 240826 162454
rect 241382 162218 280826 162454
rect 281382 162218 320826 162454
rect 321062 162218 321146 162454
rect 321382 162218 360826 162454
rect 361062 162218 361146 162454
rect 361382 162218 400826 162454
rect 401062 162218 401146 162454
rect 401382 162218 440826 162454
rect 441062 162218 441146 162454
rect 441382 162218 480826 162454
rect 481062 162218 481146 162454
rect 481382 162218 520826 162454
rect 521062 162218 521146 162454
rect 521382 162218 560826 162454
rect 561062 162218 561146 162454
rect 561382 162218 585342 162454
rect 585578 162218 585662 162454
rect 585898 162218 586890 162454
rect -2966 162134 586890 162218
rect -2966 161898 -1974 162134
rect -1738 161898 -1654 162134
rect -1418 161898 826 162134
rect 1062 161898 1146 162134
rect 1382 161898 40826 162134
rect 41062 161898 41146 162134
rect 41382 161898 80826 162134
rect 81062 161898 81146 162134
rect 81382 161898 120826 162134
rect 121062 161898 121146 162134
rect 121382 161898 160826 162134
rect 161382 161898 200826 162134
rect 201382 161898 240826 162134
rect 241382 161898 280826 162134
rect 281382 161898 320826 162134
rect 321062 161898 321146 162134
rect 321382 161898 360826 162134
rect 361062 161898 361146 162134
rect 361382 161898 400826 162134
rect 401062 161898 401146 162134
rect 401382 161898 440826 162134
rect 441062 161898 441146 162134
rect 441382 161898 480826 162134
rect 481062 161898 481146 162134
rect 481382 161898 520826 162134
rect 521062 161898 521146 162134
rect 521382 161898 560826 162134
rect 561062 161898 561146 162134
rect 561382 161898 585342 162134
rect 585578 161898 585662 162134
rect 585898 161898 586890 162134
rect -2966 161866 586890 161898
rect -8726 153614 592650 153646
rect -8726 153378 -8694 153614
rect -8458 153378 -8374 153614
rect -8138 153378 31986 153614
rect 32222 153378 32306 153614
rect 32542 153378 71986 153614
rect 72222 153378 72306 153614
rect 72542 153378 111986 153614
rect 112222 153378 112306 153614
rect 112542 153378 151986 153614
rect 152222 153378 152306 153614
rect 152542 153378 191986 153614
rect 192222 153378 192306 153614
rect 192542 153378 231986 153614
rect 232222 153378 232306 153614
rect 232542 153378 271986 153614
rect 272222 153378 272306 153614
rect 272542 153378 311986 153614
rect 312222 153378 312306 153614
rect 312542 153378 351986 153614
rect 352222 153378 352306 153614
rect 352542 153378 391986 153614
rect 392222 153378 392306 153614
rect 392542 153378 431986 153614
rect 432222 153378 432306 153614
rect 432542 153378 471986 153614
rect 472222 153378 472306 153614
rect 472542 153378 511986 153614
rect 512222 153378 512306 153614
rect 512542 153378 551986 153614
rect 552222 153378 552306 153614
rect 552542 153378 592062 153614
rect 592298 153378 592382 153614
rect 592618 153378 592650 153614
rect -8726 153294 592650 153378
rect -8726 153058 -8694 153294
rect -8458 153058 -8374 153294
rect -8138 153058 31986 153294
rect 32222 153058 32306 153294
rect 32542 153058 71986 153294
rect 72222 153058 72306 153294
rect 72542 153058 111986 153294
rect 112222 153058 112306 153294
rect 112542 153058 151986 153294
rect 152222 153058 152306 153294
rect 152542 153058 191986 153294
rect 192222 153058 192306 153294
rect 192542 153058 231986 153294
rect 232222 153058 232306 153294
rect 232542 153058 271986 153294
rect 272222 153058 272306 153294
rect 272542 153058 311986 153294
rect 312222 153058 312306 153294
rect 312542 153058 351986 153294
rect 352222 153058 352306 153294
rect 352542 153058 391986 153294
rect 392222 153058 392306 153294
rect 392542 153058 431986 153294
rect 432222 153058 432306 153294
rect 432542 153058 471986 153294
rect 472222 153058 472306 153294
rect 472542 153058 511986 153294
rect 512222 153058 512306 153294
rect 512542 153058 551986 153294
rect 552222 153058 552306 153294
rect 552542 153058 592062 153294
rect 592298 153058 592382 153294
rect 592618 153058 592650 153294
rect -8726 153026 592650 153058
rect -6806 149894 590730 149926
rect -6806 149658 -6774 149894
rect -6538 149658 -6454 149894
rect -6218 149658 28266 149894
rect 28502 149658 28586 149894
rect 28822 149658 68266 149894
rect 68502 149658 68586 149894
rect 68822 149658 108266 149894
rect 108502 149658 108586 149894
rect 108822 149658 148266 149894
rect 148502 149658 148586 149894
rect 148822 149658 188266 149894
rect 188502 149658 188586 149894
rect 188822 149658 228266 149894
rect 228502 149658 228586 149894
rect 228822 149658 268266 149894
rect 268502 149658 268586 149894
rect 268822 149658 308266 149894
rect 308502 149658 308586 149894
rect 308822 149658 348266 149894
rect 348502 149658 348586 149894
rect 348822 149658 388266 149894
rect 388502 149658 388586 149894
rect 388822 149658 428266 149894
rect 428502 149658 428586 149894
rect 428822 149658 468266 149894
rect 468502 149658 468586 149894
rect 468822 149658 508266 149894
rect 508502 149658 508586 149894
rect 508822 149658 548266 149894
rect 548502 149658 548586 149894
rect 548822 149658 590142 149894
rect 590378 149658 590462 149894
rect 590698 149658 590730 149894
rect -6806 149574 590730 149658
rect -6806 149338 -6774 149574
rect -6538 149338 -6454 149574
rect -6218 149338 28266 149574
rect 28502 149338 28586 149574
rect 28822 149338 68266 149574
rect 68502 149338 68586 149574
rect 68822 149338 108266 149574
rect 108502 149338 108586 149574
rect 108822 149338 148266 149574
rect 148502 149338 148586 149574
rect 148822 149338 188266 149574
rect 188502 149338 188586 149574
rect 188822 149338 228266 149574
rect 228502 149338 228586 149574
rect 228822 149338 268266 149574
rect 268502 149338 268586 149574
rect 268822 149338 308266 149574
rect 308502 149338 308586 149574
rect 308822 149338 348266 149574
rect 348502 149338 348586 149574
rect 348822 149338 388266 149574
rect 388502 149338 388586 149574
rect 388822 149338 428266 149574
rect 428502 149338 428586 149574
rect 428822 149338 468266 149574
rect 468502 149338 468586 149574
rect 468822 149338 508266 149574
rect 508502 149338 508586 149574
rect 508822 149338 548266 149574
rect 548502 149338 548586 149574
rect 548822 149338 590142 149574
rect 590378 149338 590462 149574
rect 590698 149338 590730 149574
rect -6806 149306 590730 149338
rect -4886 146174 588810 146206
rect -4886 145938 -4854 146174
rect -4618 145938 -4534 146174
rect -4298 145938 24546 146174
rect 24782 145938 24866 146174
rect 25102 145938 64546 146174
rect 64782 145938 64866 146174
rect 65102 145938 104546 146174
rect 104782 145938 104866 146174
rect 105102 145938 144546 146174
rect 144782 145938 144866 146174
rect 145102 145938 184546 146174
rect 184782 145938 184866 146174
rect 185102 145938 224546 146174
rect 224782 145938 224866 146174
rect 225102 145938 264546 146174
rect 264782 145938 264866 146174
rect 265102 145938 304546 146174
rect 304782 145938 304866 146174
rect 305102 145938 344546 146174
rect 344782 145938 344866 146174
rect 345102 145938 384546 146174
rect 384782 145938 384866 146174
rect 385102 145938 424546 146174
rect 424782 145938 424866 146174
rect 425102 145938 464546 146174
rect 464782 145938 464866 146174
rect 465102 145938 504546 146174
rect 504782 145938 504866 146174
rect 505102 145938 544546 146174
rect 544782 145938 544866 146174
rect 545102 145938 588222 146174
rect 588458 145938 588542 146174
rect 588778 145938 588810 146174
rect -4886 145854 588810 145938
rect -4886 145618 -4854 145854
rect -4618 145618 -4534 145854
rect -4298 145618 24546 145854
rect 24782 145618 24866 145854
rect 25102 145618 64546 145854
rect 64782 145618 64866 145854
rect 65102 145618 104546 145854
rect 104782 145618 104866 145854
rect 105102 145618 144546 145854
rect 144782 145618 144866 145854
rect 145102 145618 184546 145854
rect 184782 145618 184866 145854
rect 185102 145618 224546 145854
rect 224782 145618 224866 145854
rect 225102 145618 264546 145854
rect 264782 145618 264866 145854
rect 265102 145618 304546 145854
rect 304782 145618 304866 145854
rect 305102 145618 344546 145854
rect 344782 145618 344866 145854
rect 345102 145618 384546 145854
rect 384782 145618 384866 145854
rect 385102 145618 424546 145854
rect 424782 145618 424866 145854
rect 425102 145618 464546 145854
rect 464782 145618 464866 145854
rect 465102 145618 504546 145854
rect 504782 145618 504866 145854
rect 505102 145618 544546 145854
rect 544782 145618 544866 145854
rect 545102 145618 588222 145854
rect 588458 145618 588542 145854
rect 588778 145618 588810 145854
rect -4886 145586 588810 145618
rect -2966 142454 586890 142486
rect -2966 142218 -2934 142454
rect -2698 142218 -2614 142454
rect -2378 142218 20826 142454
rect 21062 142218 21146 142454
rect 21382 142218 60826 142454
rect 61062 142218 61146 142454
rect 61382 142218 100826 142454
rect 101062 142218 101146 142454
rect 101382 142218 140826 142454
rect 141382 142218 180826 142454
rect 181382 142218 220826 142454
rect 221382 142218 260826 142454
rect 261382 142218 300826 142454
rect 301382 142218 340826 142454
rect 341062 142218 341146 142454
rect 341382 142218 380826 142454
rect 381062 142218 381146 142454
rect 381382 142218 420826 142454
rect 421062 142218 421146 142454
rect 421382 142218 460826 142454
rect 461062 142218 461146 142454
rect 461382 142218 500826 142454
rect 501062 142218 501146 142454
rect 501382 142218 540826 142454
rect 541062 142218 541146 142454
rect 541382 142218 580826 142454
rect 581062 142218 581146 142454
rect 581382 142218 586302 142454
rect 586538 142218 586622 142454
rect 586858 142218 586890 142454
rect -2966 142134 586890 142218
rect -2966 141898 -2934 142134
rect -2698 141898 -2614 142134
rect -2378 141898 20826 142134
rect 21062 141898 21146 142134
rect 21382 141898 60826 142134
rect 61062 141898 61146 142134
rect 61382 141898 100826 142134
rect 101062 141898 101146 142134
rect 101382 141898 140826 142134
rect 141382 141898 180826 142134
rect 181382 141898 220826 142134
rect 221382 141898 260826 142134
rect 261382 141898 300826 142134
rect 301382 141898 340826 142134
rect 341062 141898 341146 142134
rect 341382 141898 380826 142134
rect 381062 141898 381146 142134
rect 381382 141898 420826 142134
rect 421062 141898 421146 142134
rect 421382 141898 460826 142134
rect 461062 141898 461146 142134
rect 461382 141898 500826 142134
rect 501062 141898 501146 142134
rect 501382 141898 540826 142134
rect 541062 141898 541146 142134
rect 541382 141898 580826 142134
rect 581062 141898 581146 142134
rect 581382 141898 586302 142134
rect 586538 141898 586622 142134
rect 586858 141898 586890 142134
rect -2966 141866 586890 141898
rect -8726 133614 592650 133646
rect -8726 133378 -7734 133614
rect -7498 133378 -7414 133614
rect -7178 133378 11986 133614
rect 12222 133378 12306 133614
rect 12542 133378 51986 133614
rect 52222 133378 52306 133614
rect 52542 133378 91986 133614
rect 92222 133378 92306 133614
rect 92542 133378 131986 133614
rect 132222 133378 132306 133614
rect 132542 133378 171986 133614
rect 172222 133378 172306 133614
rect 172542 133378 211986 133614
rect 212222 133378 212306 133614
rect 212542 133378 251986 133614
rect 252222 133378 252306 133614
rect 252542 133378 291986 133614
rect 292222 133378 292306 133614
rect 292542 133378 331986 133614
rect 332222 133378 332306 133614
rect 332542 133378 371986 133614
rect 372222 133378 372306 133614
rect 372542 133378 411986 133614
rect 412222 133378 412306 133614
rect 412542 133378 451986 133614
rect 452222 133378 452306 133614
rect 452542 133378 491986 133614
rect 492222 133378 492306 133614
rect 492542 133378 531986 133614
rect 532222 133378 532306 133614
rect 532542 133378 571986 133614
rect 572222 133378 572306 133614
rect 572542 133378 591102 133614
rect 591338 133378 591422 133614
rect 591658 133378 592650 133614
rect -8726 133294 592650 133378
rect -8726 133058 -7734 133294
rect -7498 133058 -7414 133294
rect -7178 133058 11986 133294
rect 12222 133058 12306 133294
rect 12542 133058 51986 133294
rect 52222 133058 52306 133294
rect 52542 133058 91986 133294
rect 92222 133058 92306 133294
rect 92542 133058 131986 133294
rect 132222 133058 132306 133294
rect 132542 133058 171986 133294
rect 172222 133058 172306 133294
rect 172542 133058 211986 133294
rect 212222 133058 212306 133294
rect 212542 133058 251986 133294
rect 252222 133058 252306 133294
rect 252542 133058 291986 133294
rect 292222 133058 292306 133294
rect 292542 133058 331986 133294
rect 332222 133058 332306 133294
rect 332542 133058 371986 133294
rect 372222 133058 372306 133294
rect 372542 133058 411986 133294
rect 412222 133058 412306 133294
rect 412542 133058 451986 133294
rect 452222 133058 452306 133294
rect 452542 133058 491986 133294
rect 492222 133058 492306 133294
rect 492542 133058 531986 133294
rect 532222 133058 532306 133294
rect 532542 133058 571986 133294
rect 572222 133058 572306 133294
rect 572542 133058 591102 133294
rect 591338 133058 591422 133294
rect 591658 133058 592650 133294
rect -8726 133026 592650 133058
rect -6806 129894 590730 129926
rect -6806 129658 -5814 129894
rect -5578 129658 -5494 129894
rect -5258 129658 8266 129894
rect 8502 129658 8586 129894
rect 8822 129658 48266 129894
rect 48502 129658 48586 129894
rect 48822 129658 88266 129894
rect 88502 129658 88586 129894
rect 88822 129658 128266 129894
rect 128502 129658 128586 129894
rect 128822 129658 168266 129894
rect 168502 129658 168586 129894
rect 168822 129658 208266 129894
rect 208502 129658 208586 129894
rect 208822 129658 248266 129894
rect 248502 129658 248586 129894
rect 248822 129658 288266 129894
rect 288502 129658 288586 129894
rect 288822 129658 328266 129894
rect 328502 129658 328586 129894
rect 328822 129658 368266 129894
rect 368502 129658 368586 129894
rect 368822 129658 408266 129894
rect 408502 129658 408586 129894
rect 408822 129658 448266 129894
rect 448502 129658 448586 129894
rect 448822 129658 488266 129894
rect 488502 129658 488586 129894
rect 488822 129658 528266 129894
rect 528502 129658 528586 129894
rect 528822 129658 568266 129894
rect 568502 129658 568586 129894
rect 568822 129658 589182 129894
rect 589418 129658 589502 129894
rect 589738 129658 590730 129894
rect -6806 129574 590730 129658
rect -6806 129338 -5814 129574
rect -5578 129338 -5494 129574
rect -5258 129338 8266 129574
rect 8502 129338 8586 129574
rect 8822 129338 48266 129574
rect 48502 129338 48586 129574
rect 48822 129338 88266 129574
rect 88502 129338 88586 129574
rect 88822 129338 128266 129574
rect 128502 129338 128586 129574
rect 128822 129338 168266 129574
rect 168502 129338 168586 129574
rect 168822 129338 208266 129574
rect 208502 129338 208586 129574
rect 208822 129338 248266 129574
rect 248502 129338 248586 129574
rect 248822 129338 288266 129574
rect 288502 129338 288586 129574
rect 288822 129338 328266 129574
rect 328502 129338 328586 129574
rect 328822 129338 368266 129574
rect 368502 129338 368586 129574
rect 368822 129338 408266 129574
rect 408502 129338 408586 129574
rect 408822 129338 448266 129574
rect 448502 129338 448586 129574
rect 448822 129338 488266 129574
rect 488502 129338 488586 129574
rect 488822 129338 528266 129574
rect 528502 129338 528586 129574
rect 528822 129338 568266 129574
rect 568502 129338 568586 129574
rect 568822 129338 589182 129574
rect 589418 129338 589502 129574
rect 589738 129338 590730 129574
rect -6806 129306 590730 129338
rect -4886 126174 588810 126206
rect -4886 125938 -3894 126174
rect -3658 125938 -3574 126174
rect -3338 125938 4546 126174
rect 4782 125938 4866 126174
rect 5102 125938 44546 126174
rect 44782 125938 44866 126174
rect 45102 125938 84546 126174
rect 84782 125938 84866 126174
rect 85102 125938 124546 126174
rect 124782 125938 124866 126174
rect 125102 125938 164546 126174
rect 164782 125938 164866 126174
rect 165102 125938 204546 126174
rect 204782 125938 204866 126174
rect 205102 125938 244546 126174
rect 244782 125938 244866 126174
rect 245102 125938 284546 126174
rect 284782 125938 284866 126174
rect 285102 125938 324546 126174
rect 324782 125938 324866 126174
rect 325102 125938 364546 126174
rect 364782 125938 364866 126174
rect 365102 125938 404546 126174
rect 404782 125938 404866 126174
rect 405102 125938 444546 126174
rect 444782 125938 444866 126174
rect 445102 125938 484546 126174
rect 484782 125938 484866 126174
rect 485102 125938 524546 126174
rect 524782 125938 524866 126174
rect 525102 125938 564546 126174
rect 564782 125938 564866 126174
rect 565102 125938 587262 126174
rect 587498 125938 587582 126174
rect 587818 125938 588810 126174
rect -4886 125854 588810 125938
rect -4886 125618 -3894 125854
rect -3658 125618 -3574 125854
rect -3338 125618 4546 125854
rect 4782 125618 4866 125854
rect 5102 125618 44546 125854
rect 44782 125618 44866 125854
rect 45102 125618 84546 125854
rect 84782 125618 84866 125854
rect 85102 125618 124546 125854
rect 124782 125618 124866 125854
rect 125102 125618 164546 125854
rect 164782 125618 164866 125854
rect 165102 125618 204546 125854
rect 204782 125618 204866 125854
rect 205102 125618 244546 125854
rect 244782 125618 244866 125854
rect 245102 125618 284546 125854
rect 284782 125618 284866 125854
rect 285102 125618 324546 125854
rect 324782 125618 324866 125854
rect 325102 125618 364546 125854
rect 364782 125618 364866 125854
rect 365102 125618 404546 125854
rect 404782 125618 404866 125854
rect 405102 125618 444546 125854
rect 444782 125618 444866 125854
rect 445102 125618 484546 125854
rect 484782 125618 484866 125854
rect 485102 125618 524546 125854
rect 524782 125618 524866 125854
rect 525102 125618 564546 125854
rect 564782 125618 564866 125854
rect 565102 125618 587262 125854
rect 587498 125618 587582 125854
rect 587818 125618 588810 125854
rect -4886 125586 588810 125618
rect -2966 122454 586890 122486
rect -2966 122218 -1974 122454
rect -1738 122218 -1654 122454
rect -1418 122218 826 122454
rect 1062 122218 1146 122454
rect 1382 122218 40826 122454
rect 41062 122218 41146 122454
rect 41382 122218 80826 122454
rect 81062 122218 81146 122454
rect 81382 122218 120826 122454
rect 121062 122218 121146 122454
rect 121382 122218 160826 122454
rect 161062 122218 161146 122454
rect 161382 122218 200826 122454
rect 201062 122218 201146 122454
rect 201382 122218 240826 122454
rect 241062 122218 241146 122454
rect 241382 122218 280826 122454
rect 281062 122218 281146 122454
rect 281382 122218 320826 122454
rect 321062 122218 321146 122454
rect 321382 122218 360826 122454
rect 361062 122218 361146 122454
rect 361382 122218 400826 122454
rect 401062 122218 401146 122454
rect 401382 122218 440826 122454
rect 441062 122218 441146 122454
rect 441382 122218 480826 122454
rect 481062 122218 481146 122454
rect 481382 122218 520826 122454
rect 521062 122218 521146 122454
rect 521382 122218 560826 122454
rect 561062 122218 561146 122454
rect 561382 122218 585342 122454
rect 585578 122218 585662 122454
rect 585898 122218 586890 122454
rect -2966 122134 586890 122218
rect -2966 121898 -1974 122134
rect -1738 121898 -1654 122134
rect -1418 121898 826 122134
rect 1062 121898 1146 122134
rect 1382 121898 40826 122134
rect 41062 121898 41146 122134
rect 41382 121898 80826 122134
rect 81062 121898 81146 122134
rect 81382 121898 120826 122134
rect 121062 121898 121146 122134
rect 121382 121898 160826 122134
rect 161062 121898 161146 122134
rect 161382 121898 200826 122134
rect 201062 121898 201146 122134
rect 201382 121898 240826 122134
rect 241062 121898 241146 122134
rect 241382 121898 280826 122134
rect 281062 121898 281146 122134
rect 281382 121898 320826 122134
rect 321062 121898 321146 122134
rect 321382 121898 360826 122134
rect 361062 121898 361146 122134
rect 361382 121898 400826 122134
rect 401062 121898 401146 122134
rect 401382 121898 440826 122134
rect 441062 121898 441146 122134
rect 441382 121898 480826 122134
rect 481062 121898 481146 122134
rect 481382 121898 520826 122134
rect 521062 121898 521146 122134
rect 521382 121898 560826 122134
rect 561062 121898 561146 122134
rect 561382 121898 585342 122134
rect 585578 121898 585662 122134
rect 585898 121898 586890 122134
rect -2966 121866 586890 121898
rect -8726 113614 592650 113646
rect -8726 113378 -8694 113614
rect -8458 113378 -8374 113614
rect -8138 113378 31986 113614
rect 32222 113378 32306 113614
rect 32542 113378 71986 113614
rect 72222 113378 72306 113614
rect 72542 113378 111986 113614
rect 112222 113378 112306 113614
rect 112542 113378 151986 113614
rect 152222 113378 152306 113614
rect 152542 113378 191986 113614
rect 192222 113378 192306 113614
rect 192542 113378 231986 113614
rect 232222 113378 232306 113614
rect 232542 113378 271986 113614
rect 272222 113378 272306 113614
rect 272542 113378 311986 113614
rect 312222 113378 312306 113614
rect 312542 113378 351986 113614
rect 352222 113378 352306 113614
rect 352542 113378 391986 113614
rect 392222 113378 392306 113614
rect 392542 113378 431986 113614
rect 432222 113378 432306 113614
rect 432542 113378 471986 113614
rect 472222 113378 472306 113614
rect 472542 113378 511986 113614
rect 512222 113378 512306 113614
rect 512542 113378 551986 113614
rect 552222 113378 552306 113614
rect 552542 113378 592062 113614
rect 592298 113378 592382 113614
rect 592618 113378 592650 113614
rect -8726 113294 592650 113378
rect -8726 113058 -8694 113294
rect -8458 113058 -8374 113294
rect -8138 113058 31986 113294
rect 32222 113058 32306 113294
rect 32542 113058 71986 113294
rect 72222 113058 72306 113294
rect 72542 113058 111986 113294
rect 112222 113058 112306 113294
rect 112542 113058 151986 113294
rect 152222 113058 152306 113294
rect 152542 113058 191986 113294
rect 192222 113058 192306 113294
rect 192542 113058 231986 113294
rect 232222 113058 232306 113294
rect 232542 113058 271986 113294
rect 272222 113058 272306 113294
rect 272542 113058 311986 113294
rect 312222 113058 312306 113294
rect 312542 113058 351986 113294
rect 352222 113058 352306 113294
rect 352542 113058 391986 113294
rect 392222 113058 392306 113294
rect 392542 113058 431986 113294
rect 432222 113058 432306 113294
rect 432542 113058 471986 113294
rect 472222 113058 472306 113294
rect 472542 113058 511986 113294
rect 512222 113058 512306 113294
rect 512542 113058 551986 113294
rect 552222 113058 552306 113294
rect 552542 113058 592062 113294
rect 592298 113058 592382 113294
rect 592618 113058 592650 113294
rect -8726 113026 592650 113058
rect -6806 109894 590730 109926
rect -6806 109658 -6774 109894
rect -6538 109658 -6454 109894
rect -6218 109658 28266 109894
rect 28502 109658 28586 109894
rect 28822 109658 68266 109894
rect 68502 109658 68586 109894
rect 68822 109658 108266 109894
rect 108502 109658 108586 109894
rect 108822 109658 148266 109894
rect 148502 109658 148586 109894
rect 148822 109658 188266 109894
rect 188502 109658 188586 109894
rect 188822 109658 228266 109894
rect 228502 109658 228586 109894
rect 228822 109658 268266 109894
rect 268502 109658 268586 109894
rect 268822 109658 308266 109894
rect 308502 109658 308586 109894
rect 308822 109658 348266 109894
rect 348502 109658 348586 109894
rect 348822 109658 388266 109894
rect 388502 109658 388586 109894
rect 388822 109658 428266 109894
rect 428502 109658 428586 109894
rect 428822 109658 468266 109894
rect 468502 109658 468586 109894
rect 468822 109658 508266 109894
rect 508502 109658 508586 109894
rect 508822 109658 548266 109894
rect 548502 109658 548586 109894
rect 548822 109658 590142 109894
rect 590378 109658 590462 109894
rect 590698 109658 590730 109894
rect -6806 109574 590730 109658
rect -6806 109338 -6774 109574
rect -6538 109338 -6454 109574
rect -6218 109338 28266 109574
rect 28502 109338 28586 109574
rect 28822 109338 68266 109574
rect 68502 109338 68586 109574
rect 68822 109338 108266 109574
rect 108502 109338 108586 109574
rect 108822 109338 148266 109574
rect 148502 109338 148586 109574
rect 148822 109338 188266 109574
rect 188502 109338 188586 109574
rect 188822 109338 228266 109574
rect 228502 109338 228586 109574
rect 228822 109338 268266 109574
rect 268502 109338 268586 109574
rect 268822 109338 308266 109574
rect 308502 109338 308586 109574
rect 308822 109338 348266 109574
rect 348502 109338 348586 109574
rect 348822 109338 388266 109574
rect 388502 109338 388586 109574
rect 388822 109338 428266 109574
rect 428502 109338 428586 109574
rect 428822 109338 468266 109574
rect 468502 109338 468586 109574
rect 468822 109338 508266 109574
rect 508502 109338 508586 109574
rect 508822 109338 548266 109574
rect 548502 109338 548586 109574
rect 548822 109338 590142 109574
rect 590378 109338 590462 109574
rect 590698 109338 590730 109574
rect -6806 109306 590730 109338
rect -4886 106174 588810 106206
rect -4886 105938 -4854 106174
rect -4618 105938 -4534 106174
rect -4298 105938 24546 106174
rect 24782 105938 24866 106174
rect 25102 105938 64546 106174
rect 64782 105938 64866 106174
rect 65102 105938 104546 106174
rect 104782 105938 104866 106174
rect 105102 105938 144546 106174
rect 144782 105938 144866 106174
rect 145102 105938 184546 106174
rect 184782 105938 184866 106174
rect 185102 105938 224546 106174
rect 224782 105938 224866 106174
rect 225102 105938 264546 106174
rect 264782 105938 264866 106174
rect 265102 105938 304546 106174
rect 304782 105938 304866 106174
rect 305102 105938 344546 106174
rect 344782 105938 344866 106174
rect 345102 105938 384546 106174
rect 384782 105938 384866 106174
rect 385102 105938 424546 106174
rect 424782 105938 424866 106174
rect 425102 105938 464546 106174
rect 464782 105938 464866 106174
rect 465102 105938 504546 106174
rect 504782 105938 504866 106174
rect 505102 105938 544546 106174
rect 544782 105938 544866 106174
rect 545102 105938 588222 106174
rect 588458 105938 588542 106174
rect 588778 105938 588810 106174
rect -4886 105854 588810 105938
rect -4886 105618 -4854 105854
rect -4618 105618 -4534 105854
rect -4298 105618 24546 105854
rect 24782 105618 24866 105854
rect 25102 105618 64546 105854
rect 64782 105618 64866 105854
rect 65102 105618 104546 105854
rect 104782 105618 104866 105854
rect 105102 105618 144546 105854
rect 144782 105618 144866 105854
rect 145102 105618 184546 105854
rect 184782 105618 184866 105854
rect 185102 105618 224546 105854
rect 224782 105618 224866 105854
rect 225102 105618 264546 105854
rect 264782 105618 264866 105854
rect 265102 105618 304546 105854
rect 304782 105618 304866 105854
rect 305102 105618 344546 105854
rect 344782 105618 344866 105854
rect 345102 105618 384546 105854
rect 384782 105618 384866 105854
rect 385102 105618 424546 105854
rect 424782 105618 424866 105854
rect 425102 105618 464546 105854
rect 464782 105618 464866 105854
rect 465102 105618 504546 105854
rect 504782 105618 504866 105854
rect 505102 105618 544546 105854
rect 544782 105618 544866 105854
rect 545102 105618 588222 105854
rect 588458 105618 588542 105854
rect 588778 105618 588810 105854
rect -4886 105586 588810 105618
rect -2966 102454 586890 102486
rect -2966 102218 -2934 102454
rect -2698 102218 -2614 102454
rect -2378 102218 20826 102454
rect 21062 102218 21146 102454
rect 21382 102218 60826 102454
rect 61062 102218 61146 102454
rect 61382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 140826 102454
rect 141062 102218 141146 102454
rect 141382 102218 180826 102454
rect 181062 102218 181146 102454
rect 181382 102218 220826 102454
rect 221062 102218 221146 102454
rect 221382 102218 260826 102454
rect 261062 102218 261146 102454
rect 261382 102218 300826 102454
rect 301062 102218 301146 102454
rect 301382 102218 340826 102454
rect 341062 102218 341146 102454
rect 341382 102218 380826 102454
rect 381062 102218 381146 102454
rect 381382 102218 420826 102454
rect 421062 102218 421146 102454
rect 421382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 500826 102454
rect 501062 102218 501146 102454
rect 501382 102218 540826 102454
rect 541062 102218 541146 102454
rect 541382 102218 580826 102454
rect 581062 102218 581146 102454
rect 581382 102218 586302 102454
rect 586538 102218 586622 102454
rect 586858 102218 586890 102454
rect -2966 102134 586890 102218
rect -2966 101898 -2934 102134
rect -2698 101898 -2614 102134
rect -2378 101898 20826 102134
rect 21062 101898 21146 102134
rect 21382 101898 60826 102134
rect 61062 101898 61146 102134
rect 61382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 140826 102134
rect 141062 101898 141146 102134
rect 141382 101898 180826 102134
rect 181062 101898 181146 102134
rect 181382 101898 220826 102134
rect 221062 101898 221146 102134
rect 221382 101898 260826 102134
rect 261062 101898 261146 102134
rect 261382 101898 300826 102134
rect 301062 101898 301146 102134
rect 301382 101898 340826 102134
rect 341062 101898 341146 102134
rect 341382 101898 380826 102134
rect 381062 101898 381146 102134
rect 381382 101898 420826 102134
rect 421062 101898 421146 102134
rect 421382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 500826 102134
rect 501062 101898 501146 102134
rect 501382 101898 540826 102134
rect 541062 101898 541146 102134
rect 541382 101898 580826 102134
rect 581062 101898 581146 102134
rect 581382 101898 586302 102134
rect 586538 101898 586622 102134
rect 586858 101898 586890 102134
rect -2966 101866 586890 101898
rect -8726 93614 592650 93646
rect -8726 93378 -7734 93614
rect -7498 93378 -7414 93614
rect -7178 93378 11986 93614
rect 12222 93378 12306 93614
rect 12542 93378 51986 93614
rect 52222 93378 52306 93614
rect 52542 93378 91986 93614
rect 92222 93378 92306 93614
rect 92542 93378 131986 93614
rect 132222 93378 132306 93614
rect 132542 93378 171986 93614
rect 172222 93378 172306 93614
rect 172542 93378 211986 93614
rect 212222 93378 212306 93614
rect 212542 93378 251986 93614
rect 252222 93378 252306 93614
rect 252542 93378 291986 93614
rect 292222 93378 292306 93614
rect 292542 93378 331986 93614
rect 332222 93378 332306 93614
rect 332542 93378 371986 93614
rect 372222 93378 372306 93614
rect 372542 93378 411986 93614
rect 412222 93378 412306 93614
rect 412542 93378 451986 93614
rect 452222 93378 452306 93614
rect 452542 93378 491986 93614
rect 492222 93378 492306 93614
rect 492542 93378 531986 93614
rect 532222 93378 532306 93614
rect 532542 93378 571986 93614
rect 572222 93378 572306 93614
rect 572542 93378 591102 93614
rect 591338 93378 591422 93614
rect 591658 93378 592650 93614
rect -8726 93294 592650 93378
rect -8726 93058 -7734 93294
rect -7498 93058 -7414 93294
rect -7178 93058 11986 93294
rect 12222 93058 12306 93294
rect 12542 93058 51986 93294
rect 52222 93058 52306 93294
rect 52542 93058 91986 93294
rect 92222 93058 92306 93294
rect 92542 93058 131986 93294
rect 132222 93058 132306 93294
rect 132542 93058 171986 93294
rect 172222 93058 172306 93294
rect 172542 93058 211986 93294
rect 212222 93058 212306 93294
rect 212542 93058 251986 93294
rect 252222 93058 252306 93294
rect 252542 93058 291986 93294
rect 292222 93058 292306 93294
rect 292542 93058 331986 93294
rect 332222 93058 332306 93294
rect 332542 93058 371986 93294
rect 372222 93058 372306 93294
rect 372542 93058 411986 93294
rect 412222 93058 412306 93294
rect 412542 93058 451986 93294
rect 452222 93058 452306 93294
rect 452542 93058 491986 93294
rect 492222 93058 492306 93294
rect 492542 93058 531986 93294
rect 532222 93058 532306 93294
rect 532542 93058 571986 93294
rect 572222 93058 572306 93294
rect 572542 93058 591102 93294
rect 591338 93058 591422 93294
rect 591658 93058 592650 93294
rect -8726 93026 592650 93058
rect -6806 89894 590730 89926
rect -6806 89658 -5814 89894
rect -5578 89658 -5494 89894
rect -5258 89658 8266 89894
rect 8502 89658 8586 89894
rect 8822 89658 48266 89894
rect 48502 89658 48586 89894
rect 48822 89658 88266 89894
rect 88502 89658 88586 89894
rect 88822 89658 128266 89894
rect 128502 89658 128586 89894
rect 128822 89658 168266 89894
rect 168502 89658 168586 89894
rect 168822 89658 208266 89894
rect 208502 89658 208586 89894
rect 208822 89658 248266 89894
rect 248502 89658 248586 89894
rect 248822 89658 288266 89894
rect 288502 89658 288586 89894
rect 288822 89658 328266 89894
rect 328502 89658 328586 89894
rect 328822 89658 368266 89894
rect 368502 89658 368586 89894
rect 368822 89658 408266 89894
rect 408502 89658 408586 89894
rect 408822 89658 448266 89894
rect 448502 89658 448586 89894
rect 448822 89658 488266 89894
rect 488502 89658 488586 89894
rect 488822 89658 528266 89894
rect 528502 89658 528586 89894
rect 528822 89658 568266 89894
rect 568502 89658 568586 89894
rect 568822 89658 589182 89894
rect 589418 89658 589502 89894
rect 589738 89658 590730 89894
rect -6806 89574 590730 89658
rect -6806 89338 -5814 89574
rect -5578 89338 -5494 89574
rect -5258 89338 8266 89574
rect 8502 89338 8586 89574
rect 8822 89338 48266 89574
rect 48502 89338 48586 89574
rect 48822 89338 88266 89574
rect 88502 89338 88586 89574
rect 88822 89338 128266 89574
rect 128502 89338 128586 89574
rect 128822 89338 168266 89574
rect 168502 89338 168586 89574
rect 168822 89338 208266 89574
rect 208502 89338 208586 89574
rect 208822 89338 248266 89574
rect 248502 89338 248586 89574
rect 248822 89338 288266 89574
rect 288502 89338 288586 89574
rect 288822 89338 328266 89574
rect 328502 89338 328586 89574
rect 328822 89338 368266 89574
rect 368502 89338 368586 89574
rect 368822 89338 408266 89574
rect 408502 89338 408586 89574
rect 408822 89338 448266 89574
rect 448502 89338 448586 89574
rect 448822 89338 488266 89574
rect 488502 89338 488586 89574
rect 488822 89338 528266 89574
rect 528502 89338 528586 89574
rect 528822 89338 568266 89574
rect 568502 89338 568586 89574
rect 568822 89338 589182 89574
rect 589418 89338 589502 89574
rect 589738 89338 590730 89574
rect -6806 89306 590730 89338
rect -4886 86174 588810 86206
rect -4886 85938 -3894 86174
rect -3658 85938 -3574 86174
rect -3338 85938 4546 86174
rect 4782 85938 4866 86174
rect 5102 85938 44546 86174
rect 44782 85938 44866 86174
rect 45102 85938 84546 86174
rect 84782 85938 84866 86174
rect 85102 85938 124546 86174
rect 124782 85938 124866 86174
rect 125102 85938 164546 86174
rect 164782 85938 164866 86174
rect 165102 85938 204546 86174
rect 204782 85938 204866 86174
rect 205102 85938 244546 86174
rect 244782 85938 244866 86174
rect 245102 85938 284546 86174
rect 284782 85938 284866 86174
rect 285102 85938 324546 86174
rect 324782 85938 324866 86174
rect 325102 85938 364546 86174
rect 364782 85938 364866 86174
rect 365102 85938 404546 86174
rect 404782 85938 404866 86174
rect 405102 85938 444546 86174
rect 444782 85938 444866 86174
rect 445102 85938 484546 86174
rect 484782 85938 484866 86174
rect 485102 85938 524546 86174
rect 524782 85938 524866 86174
rect 525102 85938 564546 86174
rect 564782 85938 564866 86174
rect 565102 85938 587262 86174
rect 587498 85938 587582 86174
rect 587818 85938 588810 86174
rect -4886 85854 588810 85938
rect -4886 85618 -3894 85854
rect -3658 85618 -3574 85854
rect -3338 85618 4546 85854
rect 4782 85618 4866 85854
rect 5102 85618 44546 85854
rect 44782 85618 44866 85854
rect 45102 85618 84546 85854
rect 84782 85618 84866 85854
rect 85102 85618 124546 85854
rect 124782 85618 124866 85854
rect 125102 85618 164546 85854
rect 164782 85618 164866 85854
rect 165102 85618 204546 85854
rect 204782 85618 204866 85854
rect 205102 85618 244546 85854
rect 244782 85618 244866 85854
rect 245102 85618 284546 85854
rect 284782 85618 284866 85854
rect 285102 85618 324546 85854
rect 324782 85618 324866 85854
rect 325102 85618 364546 85854
rect 364782 85618 364866 85854
rect 365102 85618 404546 85854
rect 404782 85618 404866 85854
rect 405102 85618 444546 85854
rect 444782 85618 444866 85854
rect 445102 85618 484546 85854
rect 484782 85618 484866 85854
rect 485102 85618 524546 85854
rect 524782 85618 524866 85854
rect 525102 85618 564546 85854
rect 564782 85618 564866 85854
rect 565102 85618 587262 85854
rect 587498 85618 587582 85854
rect 587818 85618 588810 85854
rect -4886 85586 588810 85618
rect -2966 82454 586890 82486
rect -2966 82218 -1974 82454
rect -1738 82218 -1654 82454
rect -1418 82218 826 82454
rect 1062 82218 1146 82454
rect 1382 82218 40826 82454
rect 41062 82218 41146 82454
rect 41382 82218 80826 82454
rect 81062 82218 81146 82454
rect 81382 82218 120826 82454
rect 121062 82218 121146 82454
rect 121382 82218 160826 82454
rect 161062 82218 161146 82454
rect 161382 82218 200826 82454
rect 201062 82218 201146 82454
rect 201382 82218 240826 82454
rect 241062 82218 241146 82454
rect 241382 82218 280826 82454
rect 281062 82218 281146 82454
rect 281382 82218 320826 82454
rect 321062 82218 321146 82454
rect 321382 82218 360826 82454
rect 361062 82218 361146 82454
rect 361382 82218 400826 82454
rect 401062 82218 401146 82454
rect 401382 82218 440826 82454
rect 441062 82218 441146 82454
rect 441382 82218 480826 82454
rect 481062 82218 481146 82454
rect 481382 82218 520826 82454
rect 521062 82218 521146 82454
rect 521382 82218 560826 82454
rect 561062 82218 561146 82454
rect 561382 82218 585342 82454
rect 585578 82218 585662 82454
rect 585898 82218 586890 82454
rect -2966 82134 586890 82218
rect -2966 81898 -1974 82134
rect -1738 81898 -1654 82134
rect -1418 81898 826 82134
rect 1062 81898 1146 82134
rect 1382 81898 40826 82134
rect 41062 81898 41146 82134
rect 41382 81898 80826 82134
rect 81062 81898 81146 82134
rect 81382 81898 120826 82134
rect 121062 81898 121146 82134
rect 121382 81898 160826 82134
rect 161062 81898 161146 82134
rect 161382 81898 200826 82134
rect 201062 81898 201146 82134
rect 201382 81898 240826 82134
rect 241062 81898 241146 82134
rect 241382 81898 280826 82134
rect 281062 81898 281146 82134
rect 281382 81898 320826 82134
rect 321062 81898 321146 82134
rect 321382 81898 360826 82134
rect 361062 81898 361146 82134
rect 361382 81898 400826 82134
rect 401062 81898 401146 82134
rect 401382 81898 440826 82134
rect 441062 81898 441146 82134
rect 441382 81898 480826 82134
rect 481062 81898 481146 82134
rect 481382 81898 520826 82134
rect 521062 81898 521146 82134
rect 521382 81898 560826 82134
rect 561062 81898 561146 82134
rect 561382 81898 585342 82134
rect 585578 81898 585662 82134
rect 585898 81898 586890 82134
rect -2966 81866 586890 81898
rect -8726 73614 592650 73646
rect -8726 73378 -8694 73614
rect -8458 73378 -8374 73614
rect -8138 73378 31986 73614
rect 32222 73378 32306 73614
rect 32542 73378 71986 73614
rect 72222 73378 72306 73614
rect 72542 73378 111986 73614
rect 112222 73378 112306 73614
rect 112542 73378 151986 73614
rect 152222 73378 152306 73614
rect 152542 73378 191986 73614
rect 192222 73378 192306 73614
rect 192542 73378 231986 73614
rect 232222 73378 232306 73614
rect 232542 73378 271986 73614
rect 272222 73378 272306 73614
rect 272542 73378 311986 73614
rect 312222 73378 312306 73614
rect 312542 73378 351986 73614
rect 352222 73378 352306 73614
rect 352542 73378 391986 73614
rect 392222 73378 392306 73614
rect 392542 73378 431986 73614
rect 432222 73378 432306 73614
rect 432542 73378 471986 73614
rect 472222 73378 472306 73614
rect 472542 73378 511986 73614
rect 512222 73378 512306 73614
rect 512542 73378 551986 73614
rect 552222 73378 552306 73614
rect 552542 73378 592062 73614
rect 592298 73378 592382 73614
rect 592618 73378 592650 73614
rect -8726 73294 592650 73378
rect -8726 73058 -8694 73294
rect -8458 73058 -8374 73294
rect -8138 73058 31986 73294
rect 32222 73058 32306 73294
rect 32542 73058 71986 73294
rect 72222 73058 72306 73294
rect 72542 73058 111986 73294
rect 112222 73058 112306 73294
rect 112542 73058 151986 73294
rect 152222 73058 152306 73294
rect 152542 73058 191986 73294
rect 192222 73058 192306 73294
rect 192542 73058 231986 73294
rect 232222 73058 232306 73294
rect 232542 73058 271986 73294
rect 272222 73058 272306 73294
rect 272542 73058 311986 73294
rect 312222 73058 312306 73294
rect 312542 73058 351986 73294
rect 352222 73058 352306 73294
rect 352542 73058 391986 73294
rect 392222 73058 392306 73294
rect 392542 73058 431986 73294
rect 432222 73058 432306 73294
rect 432542 73058 471986 73294
rect 472222 73058 472306 73294
rect 472542 73058 511986 73294
rect 512222 73058 512306 73294
rect 512542 73058 551986 73294
rect 552222 73058 552306 73294
rect 552542 73058 592062 73294
rect 592298 73058 592382 73294
rect 592618 73058 592650 73294
rect -8726 73026 592650 73058
rect -6806 69894 590730 69926
rect -6806 69658 -6774 69894
rect -6538 69658 -6454 69894
rect -6218 69658 28266 69894
rect 28502 69658 28586 69894
rect 28822 69658 68266 69894
rect 68502 69658 68586 69894
rect 68822 69658 108266 69894
rect 108502 69658 108586 69894
rect 108822 69658 148266 69894
rect 148502 69658 148586 69894
rect 148822 69658 188266 69894
rect 188502 69658 188586 69894
rect 188822 69658 228266 69894
rect 228502 69658 228586 69894
rect 228822 69658 268266 69894
rect 268502 69658 268586 69894
rect 268822 69658 308266 69894
rect 308502 69658 308586 69894
rect 308822 69658 348266 69894
rect 348502 69658 348586 69894
rect 348822 69658 388266 69894
rect 388502 69658 388586 69894
rect 388822 69658 428266 69894
rect 428502 69658 428586 69894
rect 428822 69658 468266 69894
rect 468502 69658 468586 69894
rect 468822 69658 508266 69894
rect 508502 69658 508586 69894
rect 508822 69658 548266 69894
rect 548502 69658 548586 69894
rect 548822 69658 590142 69894
rect 590378 69658 590462 69894
rect 590698 69658 590730 69894
rect -6806 69574 590730 69658
rect -6806 69338 -6774 69574
rect -6538 69338 -6454 69574
rect -6218 69338 28266 69574
rect 28502 69338 28586 69574
rect 28822 69338 68266 69574
rect 68502 69338 68586 69574
rect 68822 69338 108266 69574
rect 108502 69338 108586 69574
rect 108822 69338 148266 69574
rect 148502 69338 148586 69574
rect 148822 69338 188266 69574
rect 188502 69338 188586 69574
rect 188822 69338 228266 69574
rect 228502 69338 228586 69574
rect 228822 69338 268266 69574
rect 268502 69338 268586 69574
rect 268822 69338 308266 69574
rect 308502 69338 308586 69574
rect 308822 69338 348266 69574
rect 348502 69338 348586 69574
rect 348822 69338 388266 69574
rect 388502 69338 388586 69574
rect 388822 69338 428266 69574
rect 428502 69338 428586 69574
rect 428822 69338 468266 69574
rect 468502 69338 468586 69574
rect 468822 69338 508266 69574
rect 508502 69338 508586 69574
rect 508822 69338 548266 69574
rect 548502 69338 548586 69574
rect 548822 69338 590142 69574
rect 590378 69338 590462 69574
rect 590698 69338 590730 69574
rect -6806 69306 590730 69338
rect -4886 66174 588810 66206
rect -4886 65938 -4854 66174
rect -4618 65938 -4534 66174
rect -4298 65938 24546 66174
rect 24782 65938 24866 66174
rect 25102 65938 64546 66174
rect 64782 65938 64866 66174
rect 65102 65938 104546 66174
rect 104782 65938 104866 66174
rect 105102 65938 144546 66174
rect 144782 65938 144866 66174
rect 145102 65938 184546 66174
rect 184782 65938 184866 66174
rect 185102 65938 224546 66174
rect 224782 65938 224866 66174
rect 225102 65938 264546 66174
rect 264782 65938 264866 66174
rect 265102 65938 304546 66174
rect 304782 65938 304866 66174
rect 305102 65938 344546 66174
rect 344782 65938 344866 66174
rect 345102 65938 384546 66174
rect 384782 65938 384866 66174
rect 385102 65938 424546 66174
rect 424782 65938 424866 66174
rect 425102 65938 464546 66174
rect 464782 65938 464866 66174
rect 465102 65938 504546 66174
rect 504782 65938 504866 66174
rect 505102 65938 544546 66174
rect 544782 65938 544866 66174
rect 545102 65938 588222 66174
rect 588458 65938 588542 66174
rect 588778 65938 588810 66174
rect -4886 65854 588810 65938
rect -4886 65618 -4854 65854
rect -4618 65618 -4534 65854
rect -4298 65618 24546 65854
rect 24782 65618 24866 65854
rect 25102 65618 64546 65854
rect 64782 65618 64866 65854
rect 65102 65618 104546 65854
rect 104782 65618 104866 65854
rect 105102 65618 144546 65854
rect 144782 65618 144866 65854
rect 145102 65618 184546 65854
rect 184782 65618 184866 65854
rect 185102 65618 224546 65854
rect 224782 65618 224866 65854
rect 225102 65618 264546 65854
rect 264782 65618 264866 65854
rect 265102 65618 304546 65854
rect 304782 65618 304866 65854
rect 305102 65618 344546 65854
rect 344782 65618 344866 65854
rect 345102 65618 384546 65854
rect 384782 65618 384866 65854
rect 385102 65618 424546 65854
rect 424782 65618 424866 65854
rect 425102 65618 464546 65854
rect 464782 65618 464866 65854
rect 465102 65618 504546 65854
rect 504782 65618 504866 65854
rect 505102 65618 544546 65854
rect 544782 65618 544866 65854
rect 545102 65618 588222 65854
rect 588458 65618 588542 65854
rect 588778 65618 588810 65854
rect -4886 65586 588810 65618
rect -2966 62454 586890 62486
rect -2966 62218 -2934 62454
rect -2698 62218 -2614 62454
rect -2378 62218 20826 62454
rect 21062 62218 21146 62454
rect 21382 62218 60826 62454
rect 61062 62218 61146 62454
rect 61382 62218 100826 62454
rect 101062 62218 101146 62454
rect 101382 62218 140826 62454
rect 141062 62218 141146 62454
rect 141382 62218 180826 62454
rect 181062 62218 181146 62454
rect 181382 62218 220826 62454
rect 221062 62218 221146 62454
rect 221382 62218 260826 62454
rect 261062 62218 261146 62454
rect 261382 62218 300826 62454
rect 301062 62218 301146 62454
rect 301382 62218 340826 62454
rect 341062 62218 341146 62454
rect 341382 62218 380826 62454
rect 381062 62218 381146 62454
rect 381382 62218 420826 62454
rect 421062 62218 421146 62454
rect 421382 62218 460826 62454
rect 461062 62218 461146 62454
rect 461382 62218 500826 62454
rect 501062 62218 501146 62454
rect 501382 62218 540826 62454
rect 541062 62218 541146 62454
rect 541382 62218 580826 62454
rect 581062 62218 581146 62454
rect 581382 62218 586302 62454
rect 586538 62218 586622 62454
rect 586858 62218 586890 62454
rect -2966 62134 586890 62218
rect -2966 61898 -2934 62134
rect -2698 61898 -2614 62134
rect -2378 61898 20826 62134
rect 21062 61898 21146 62134
rect 21382 61898 60826 62134
rect 61062 61898 61146 62134
rect 61382 61898 100826 62134
rect 101062 61898 101146 62134
rect 101382 61898 140826 62134
rect 141062 61898 141146 62134
rect 141382 61898 180826 62134
rect 181062 61898 181146 62134
rect 181382 61898 220826 62134
rect 221062 61898 221146 62134
rect 221382 61898 260826 62134
rect 261062 61898 261146 62134
rect 261382 61898 300826 62134
rect 301062 61898 301146 62134
rect 301382 61898 340826 62134
rect 341062 61898 341146 62134
rect 341382 61898 380826 62134
rect 381062 61898 381146 62134
rect 381382 61898 420826 62134
rect 421062 61898 421146 62134
rect 421382 61898 460826 62134
rect 461062 61898 461146 62134
rect 461382 61898 500826 62134
rect 501062 61898 501146 62134
rect 501382 61898 540826 62134
rect 541062 61898 541146 62134
rect 541382 61898 580826 62134
rect 581062 61898 581146 62134
rect 581382 61898 586302 62134
rect 586538 61898 586622 62134
rect 586858 61898 586890 62134
rect -2966 61866 586890 61898
rect -8726 53614 592650 53646
rect -8726 53378 -7734 53614
rect -7498 53378 -7414 53614
rect -7178 53378 11986 53614
rect 12222 53378 12306 53614
rect 12542 53378 51986 53614
rect 52222 53378 52306 53614
rect 52542 53378 91986 53614
rect 92222 53378 92306 53614
rect 92542 53378 131986 53614
rect 132222 53378 132306 53614
rect 132542 53378 171986 53614
rect 172222 53378 172306 53614
rect 172542 53378 211986 53614
rect 212222 53378 212306 53614
rect 212542 53378 251986 53614
rect 252222 53378 252306 53614
rect 252542 53378 291986 53614
rect 292222 53378 292306 53614
rect 292542 53378 331986 53614
rect 332222 53378 332306 53614
rect 332542 53378 371986 53614
rect 372222 53378 372306 53614
rect 372542 53378 411986 53614
rect 412222 53378 412306 53614
rect 412542 53378 451986 53614
rect 452222 53378 452306 53614
rect 452542 53378 491986 53614
rect 492222 53378 492306 53614
rect 492542 53378 531986 53614
rect 532222 53378 532306 53614
rect 532542 53378 571986 53614
rect 572222 53378 572306 53614
rect 572542 53378 591102 53614
rect 591338 53378 591422 53614
rect 591658 53378 592650 53614
rect -8726 53294 592650 53378
rect -8726 53058 -7734 53294
rect -7498 53058 -7414 53294
rect -7178 53058 11986 53294
rect 12222 53058 12306 53294
rect 12542 53058 51986 53294
rect 52222 53058 52306 53294
rect 52542 53058 91986 53294
rect 92222 53058 92306 53294
rect 92542 53058 131986 53294
rect 132222 53058 132306 53294
rect 132542 53058 171986 53294
rect 172222 53058 172306 53294
rect 172542 53058 211986 53294
rect 212222 53058 212306 53294
rect 212542 53058 251986 53294
rect 252222 53058 252306 53294
rect 252542 53058 291986 53294
rect 292222 53058 292306 53294
rect 292542 53058 331986 53294
rect 332222 53058 332306 53294
rect 332542 53058 371986 53294
rect 372222 53058 372306 53294
rect 372542 53058 411986 53294
rect 412222 53058 412306 53294
rect 412542 53058 451986 53294
rect 452222 53058 452306 53294
rect 452542 53058 491986 53294
rect 492222 53058 492306 53294
rect 492542 53058 531986 53294
rect 532222 53058 532306 53294
rect 532542 53058 571986 53294
rect 572222 53058 572306 53294
rect 572542 53058 591102 53294
rect 591338 53058 591422 53294
rect 591658 53058 592650 53294
rect -8726 53026 592650 53058
rect -6806 49894 590730 49926
rect -6806 49658 -5814 49894
rect -5578 49658 -5494 49894
rect -5258 49658 8266 49894
rect 8502 49658 8586 49894
rect 8822 49658 48266 49894
rect 48502 49658 48586 49894
rect 48822 49658 88266 49894
rect 88502 49658 88586 49894
rect 88822 49658 128266 49894
rect 128502 49658 128586 49894
rect 128822 49658 168266 49894
rect 168502 49658 168586 49894
rect 168822 49658 208266 49894
rect 208502 49658 208586 49894
rect 208822 49658 248266 49894
rect 248502 49658 248586 49894
rect 248822 49658 288266 49894
rect 288502 49658 288586 49894
rect 288822 49658 328266 49894
rect 328502 49658 328586 49894
rect 328822 49658 368266 49894
rect 368502 49658 368586 49894
rect 368822 49658 408266 49894
rect 408502 49658 408586 49894
rect 408822 49658 448266 49894
rect 448502 49658 448586 49894
rect 448822 49658 488266 49894
rect 488502 49658 488586 49894
rect 488822 49658 528266 49894
rect 528502 49658 528586 49894
rect 528822 49658 568266 49894
rect 568502 49658 568586 49894
rect 568822 49658 589182 49894
rect 589418 49658 589502 49894
rect 589738 49658 590730 49894
rect -6806 49574 590730 49658
rect -6806 49338 -5814 49574
rect -5578 49338 -5494 49574
rect -5258 49338 8266 49574
rect 8502 49338 8586 49574
rect 8822 49338 48266 49574
rect 48502 49338 48586 49574
rect 48822 49338 88266 49574
rect 88502 49338 88586 49574
rect 88822 49338 128266 49574
rect 128502 49338 128586 49574
rect 128822 49338 168266 49574
rect 168502 49338 168586 49574
rect 168822 49338 208266 49574
rect 208502 49338 208586 49574
rect 208822 49338 248266 49574
rect 248502 49338 248586 49574
rect 248822 49338 288266 49574
rect 288502 49338 288586 49574
rect 288822 49338 328266 49574
rect 328502 49338 328586 49574
rect 328822 49338 368266 49574
rect 368502 49338 368586 49574
rect 368822 49338 408266 49574
rect 408502 49338 408586 49574
rect 408822 49338 448266 49574
rect 448502 49338 448586 49574
rect 448822 49338 488266 49574
rect 488502 49338 488586 49574
rect 488822 49338 528266 49574
rect 528502 49338 528586 49574
rect 528822 49338 568266 49574
rect 568502 49338 568586 49574
rect 568822 49338 589182 49574
rect 589418 49338 589502 49574
rect 589738 49338 590730 49574
rect -6806 49306 590730 49338
rect -4886 46174 588810 46206
rect -4886 45938 -3894 46174
rect -3658 45938 -3574 46174
rect -3338 45938 4546 46174
rect 4782 45938 4866 46174
rect 5102 45938 44546 46174
rect 44782 45938 44866 46174
rect 45102 45938 84546 46174
rect 84782 45938 84866 46174
rect 85102 45938 124546 46174
rect 124782 45938 124866 46174
rect 125102 45938 164546 46174
rect 164782 45938 164866 46174
rect 165102 45938 204546 46174
rect 204782 45938 204866 46174
rect 205102 45938 244546 46174
rect 244782 45938 244866 46174
rect 245102 45938 284546 46174
rect 284782 45938 284866 46174
rect 285102 45938 324546 46174
rect 324782 45938 324866 46174
rect 325102 45938 364546 46174
rect 364782 45938 364866 46174
rect 365102 45938 404546 46174
rect 404782 45938 404866 46174
rect 405102 45938 444546 46174
rect 444782 45938 444866 46174
rect 445102 45938 484546 46174
rect 484782 45938 484866 46174
rect 485102 45938 524546 46174
rect 524782 45938 524866 46174
rect 525102 45938 564546 46174
rect 564782 45938 564866 46174
rect 565102 45938 587262 46174
rect 587498 45938 587582 46174
rect 587818 45938 588810 46174
rect -4886 45854 588810 45938
rect -4886 45618 -3894 45854
rect -3658 45618 -3574 45854
rect -3338 45618 4546 45854
rect 4782 45618 4866 45854
rect 5102 45618 44546 45854
rect 44782 45618 44866 45854
rect 45102 45618 84546 45854
rect 84782 45618 84866 45854
rect 85102 45618 124546 45854
rect 124782 45618 124866 45854
rect 125102 45618 164546 45854
rect 164782 45618 164866 45854
rect 165102 45618 204546 45854
rect 204782 45618 204866 45854
rect 205102 45618 244546 45854
rect 244782 45618 244866 45854
rect 245102 45618 284546 45854
rect 284782 45618 284866 45854
rect 285102 45618 324546 45854
rect 324782 45618 324866 45854
rect 325102 45618 364546 45854
rect 364782 45618 364866 45854
rect 365102 45618 404546 45854
rect 404782 45618 404866 45854
rect 405102 45618 444546 45854
rect 444782 45618 444866 45854
rect 445102 45618 484546 45854
rect 484782 45618 484866 45854
rect 485102 45618 524546 45854
rect 524782 45618 524866 45854
rect 525102 45618 564546 45854
rect 564782 45618 564866 45854
rect 565102 45618 587262 45854
rect 587498 45618 587582 45854
rect 587818 45618 588810 45854
rect -4886 45586 588810 45618
rect -2966 42454 586890 42486
rect -2966 42218 -1974 42454
rect -1738 42218 -1654 42454
rect -1418 42218 826 42454
rect 1062 42218 1146 42454
rect 1382 42218 40826 42454
rect 41062 42218 41146 42454
rect 41382 42218 80826 42454
rect 81062 42218 81146 42454
rect 81382 42218 120826 42454
rect 121062 42218 121146 42454
rect 121382 42218 160826 42454
rect 161062 42218 161146 42454
rect 161382 42218 200826 42454
rect 201062 42218 201146 42454
rect 201382 42218 240826 42454
rect 241062 42218 241146 42454
rect 241382 42218 280826 42454
rect 281062 42218 281146 42454
rect 281382 42218 320826 42454
rect 321062 42218 321146 42454
rect 321382 42218 360826 42454
rect 361062 42218 361146 42454
rect 361382 42218 400826 42454
rect 401062 42218 401146 42454
rect 401382 42218 440826 42454
rect 441062 42218 441146 42454
rect 441382 42218 480826 42454
rect 481062 42218 481146 42454
rect 481382 42218 520826 42454
rect 521062 42218 521146 42454
rect 521382 42218 560826 42454
rect 561062 42218 561146 42454
rect 561382 42218 585342 42454
rect 585578 42218 585662 42454
rect 585898 42218 586890 42454
rect -2966 42134 586890 42218
rect -2966 41898 -1974 42134
rect -1738 41898 -1654 42134
rect -1418 41898 826 42134
rect 1062 41898 1146 42134
rect 1382 41898 40826 42134
rect 41062 41898 41146 42134
rect 41382 41898 80826 42134
rect 81062 41898 81146 42134
rect 81382 41898 120826 42134
rect 121062 41898 121146 42134
rect 121382 41898 160826 42134
rect 161062 41898 161146 42134
rect 161382 41898 200826 42134
rect 201062 41898 201146 42134
rect 201382 41898 240826 42134
rect 241062 41898 241146 42134
rect 241382 41898 280826 42134
rect 281062 41898 281146 42134
rect 281382 41898 320826 42134
rect 321062 41898 321146 42134
rect 321382 41898 360826 42134
rect 361062 41898 361146 42134
rect 361382 41898 400826 42134
rect 401062 41898 401146 42134
rect 401382 41898 440826 42134
rect 441062 41898 441146 42134
rect 441382 41898 480826 42134
rect 481062 41898 481146 42134
rect 481382 41898 520826 42134
rect 521062 41898 521146 42134
rect 521382 41898 560826 42134
rect 561062 41898 561146 42134
rect 561382 41898 585342 42134
rect 585578 41898 585662 42134
rect 585898 41898 586890 42134
rect -2966 41866 586890 41898
rect -8726 33614 592650 33646
rect -8726 33378 -8694 33614
rect -8458 33378 -8374 33614
rect -8138 33378 31986 33614
rect 32222 33378 32306 33614
rect 32542 33378 71986 33614
rect 72222 33378 72306 33614
rect 72542 33378 111986 33614
rect 112222 33378 112306 33614
rect 112542 33378 151986 33614
rect 152222 33378 152306 33614
rect 152542 33378 191986 33614
rect 192222 33378 192306 33614
rect 192542 33378 231986 33614
rect 232222 33378 232306 33614
rect 232542 33378 271986 33614
rect 272222 33378 272306 33614
rect 272542 33378 311986 33614
rect 312222 33378 312306 33614
rect 312542 33378 351986 33614
rect 352222 33378 352306 33614
rect 352542 33378 391986 33614
rect 392222 33378 392306 33614
rect 392542 33378 431986 33614
rect 432222 33378 432306 33614
rect 432542 33378 471986 33614
rect 472222 33378 472306 33614
rect 472542 33378 511986 33614
rect 512222 33378 512306 33614
rect 512542 33378 551986 33614
rect 552222 33378 552306 33614
rect 552542 33378 592062 33614
rect 592298 33378 592382 33614
rect 592618 33378 592650 33614
rect -8726 33294 592650 33378
rect -8726 33058 -8694 33294
rect -8458 33058 -8374 33294
rect -8138 33058 31986 33294
rect 32222 33058 32306 33294
rect 32542 33058 71986 33294
rect 72222 33058 72306 33294
rect 72542 33058 111986 33294
rect 112222 33058 112306 33294
rect 112542 33058 151986 33294
rect 152222 33058 152306 33294
rect 152542 33058 191986 33294
rect 192222 33058 192306 33294
rect 192542 33058 231986 33294
rect 232222 33058 232306 33294
rect 232542 33058 271986 33294
rect 272222 33058 272306 33294
rect 272542 33058 311986 33294
rect 312222 33058 312306 33294
rect 312542 33058 351986 33294
rect 352222 33058 352306 33294
rect 352542 33058 391986 33294
rect 392222 33058 392306 33294
rect 392542 33058 431986 33294
rect 432222 33058 432306 33294
rect 432542 33058 471986 33294
rect 472222 33058 472306 33294
rect 472542 33058 511986 33294
rect 512222 33058 512306 33294
rect 512542 33058 551986 33294
rect 552222 33058 552306 33294
rect 552542 33058 592062 33294
rect 592298 33058 592382 33294
rect 592618 33058 592650 33294
rect -8726 33026 592650 33058
rect -6806 29894 590730 29926
rect -6806 29658 -6774 29894
rect -6538 29658 -6454 29894
rect -6218 29658 28266 29894
rect 28502 29658 28586 29894
rect 28822 29658 68266 29894
rect 68502 29658 68586 29894
rect 68822 29658 108266 29894
rect 108502 29658 108586 29894
rect 108822 29658 148266 29894
rect 148502 29658 148586 29894
rect 148822 29658 188266 29894
rect 188502 29658 188586 29894
rect 188822 29658 228266 29894
rect 228502 29658 228586 29894
rect 228822 29658 268266 29894
rect 268502 29658 268586 29894
rect 268822 29658 308266 29894
rect 308502 29658 308586 29894
rect 308822 29658 348266 29894
rect 348502 29658 348586 29894
rect 348822 29658 388266 29894
rect 388502 29658 388586 29894
rect 388822 29658 428266 29894
rect 428502 29658 428586 29894
rect 428822 29658 468266 29894
rect 468502 29658 468586 29894
rect 468822 29658 508266 29894
rect 508502 29658 508586 29894
rect 508822 29658 548266 29894
rect 548502 29658 548586 29894
rect 548822 29658 590142 29894
rect 590378 29658 590462 29894
rect 590698 29658 590730 29894
rect -6806 29574 590730 29658
rect -6806 29338 -6774 29574
rect -6538 29338 -6454 29574
rect -6218 29338 28266 29574
rect 28502 29338 28586 29574
rect 28822 29338 68266 29574
rect 68502 29338 68586 29574
rect 68822 29338 108266 29574
rect 108502 29338 108586 29574
rect 108822 29338 148266 29574
rect 148502 29338 148586 29574
rect 148822 29338 188266 29574
rect 188502 29338 188586 29574
rect 188822 29338 228266 29574
rect 228502 29338 228586 29574
rect 228822 29338 268266 29574
rect 268502 29338 268586 29574
rect 268822 29338 308266 29574
rect 308502 29338 308586 29574
rect 308822 29338 348266 29574
rect 348502 29338 348586 29574
rect 348822 29338 388266 29574
rect 388502 29338 388586 29574
rect 388822 29338 428266 29574
rect 428502 29338 428586 29574
rect 428822 29338 468266 29574
rect 468502 29338 468586 29574
rect 468822 29338 508266 29574
rect 508502 29338 508586 29574
rect 508822 29338 548266 29574
rect 548502 29338 548586 29574
rect 548822 29338 590142 29574
rect 590378 29338 590462 29574
rect 590698 29338 590730 29574
rect -6806 29306 590730 29338
rect -4886 26174 588810 26206
rect -4886 25938 -4854 26174
rect -4618 25938 -4534 26174
rect -4298 25938 24546 26174
rect 24782 25938 24866 26174
rect 25102 25938 64546 26174
rect 64782 25938 64866 26174
rect 65102 25938 104546 26174
rect 104782 25938 104866 26174
rect 105102 25938 144546 26174
rect 144782 25938 144866 26174
rect 145102 25938 184546 26174
rect 184782 25938 184866 26174
rect 185102 25938 224546 26174
rect 224782 25938 224866 26174
rect 225102 25938 264546 26174
rect 264782 25938 264866 26174
rect 265102 25938 304546 26174
rect 304782 25938 304866 26174
rect 305102 25938 344546 26174
rect 344782 25938 344866 26174
rect 345102 25938 384546 26174
rect 384782 25938 384866 26174
rect 385102 25938 424546 26174
rect 424782 25938 424866 26174
rect 425102 25938 464546 26174
rect 464782 25938 464866 26174
rect 465102 25938 504546 26174
rect 504782 25938 504866 26174
rect 505102 25938 544546 26174
rect 544782 25938 544866 26174
rect 545102 25938 588222 26174
rect 588458 25938 588542 26174
rect 588778 25938 588810 26174
rect -4886 25854 588810 25938
rect -4886 25618 -4854 25854
rect -4618 25618 -4534 25854
rect -4298 25618 24546 25854
rect 24782 25618 24866 25854
rect 25102 25618 64546 25854
rect 64782 25618 64866 25854
rect 65102 25618 104546 25854
rect 104782 25618 104866 25854
rect 105102 25618 144546 25854
rect 144782 25618 144866 25854
rect 145102 25618 184546 25854
rect 184782 25618 184866 25854
rect 185102 25618 224546 25854
rect 224782 25618 224866 25854
rect 225102 25618 264546 25854
rect 264782 25618 264866 25854
rect 265102 25618 304546 25854
rect 304782 25618 304866 25854
rect 305102 25618 344546 25854
rect 344782 25618 344866 25854
rect 345102 25618 384546 25854
rect 384782 25618 384866 25854
rect 385102 25618 424546 25854
rect 424782 25618 424866 25854
rect 425102 25618 464546 25854
rect 464782 25618 464866 25854
rect 465102 25618 504546 25854
rect 504782 25618 504866 25854
rect 505102 25618 544546 25854
rect 544782 25618 544866 25854
rect 545102 25618 588222 25854
rect 588458 25618 588542 25854
rect 588778 25618 588810 25854
rect -4886 25586 588810 25618
rect -2966 22454 586890 22486
rect -2966 22218 -2934 22454
rect -2698 22218 -2614 22454
rect -2378 22218 20826 22454
rect 21062 22218 21146 22454
rect 21382 22218 60826 22454
rect 61062 22218 61146 22454
rect 61382 22218 100826 22454
rect 101062 22218 101146 22454
rect 101382 22218 140826 22454
rect 141062 22218 141146 22454
rect 141382 22218 180826 22454
rect 181062 22218 181146 22454
rect 181382 22218 220826 22454
rect 221062 22218 221146 22454
rect 221382 22218 260826 22454
rect 261062 22218 261146 22454
rect 261382 22218 300826 22454
rect 301062 22218 301146 22454
rect 301382 22218 340826 22454
rect 341062 22218 341146 22454
rect 341382 22218 380826 22454
rect 381062 22218 381146 22454
rect 381382 22218 420826 22454
rect 421062 22218 421146 22454
rect 421382 22218 460826 22454
rect 461062 22218 461146 22454
rect 461382 22218 500826 22454
rect 501062 22218 501146 22454
rect 501382 22218 540826 22454
rect 541062 22218 541146 22454
rect 541382 22218 580826 22454
rect 581062 22218 581146 22454
rect 581382 22218 586302 22454
rect 586538 22218 586622 22454
rect 586858 22218 586890 22454
rect -2966 22134 586890 22218
rect -2966 21898 -2934 22134
rect -2698 21898 -2614 22134
rect -2378 21898 20826 22134
rect 21062 21898 21146 22134
rect 21382 21898 60826 22134
rect 61062 21898 61146 22134
rect 61382 21898 100826 22134
rect 101062 21898 101146 22134
rect 101382 21898 140826 22134
rect 141062 21898 141146 22134
rect 141382 21898 180826 22134
rect 181062 21898 181146 22134
rect 181382 21898 220826 22134
rect 221062 21898 221146 22134
rect 221382 21898 260826 22134
rect 261062 21898 261146 22134
rect 261382 21898 300826 22134
rect 301062 21898 301146 22134
rect 301382 21898 340826 22134
rect 341062 21898 341146 22134
rect 341382 21898 380826 22134
rect 381062 21898 381146 22134
rect 381382 21898 420826 22134
rect 421062 21898 421146 22134
rect 421382 21898 460826 22134
rect 461062 21898 461146 22134
rect 461382 21898 500826 22134
rect 501062 21898 501146 22134
rect 501382 21898 540826 22134
rect 541062 21898 541146 22134
rect 541382 21898 580826 22134
rect 581062 21898 581146 22134
rect 581382 21898 586302 22134
rect 586538 21898 586622 22134
rect 586858 21898 586890 22134
rect -2966 21866 586890 21898
rect -8726 13614 592650 13646
rect -8726 13378 -7734 13614
rect -7498 13378 -7414 13614
rect -7178 13378 11986 13614
rect 12222 13378 12306 13614
rect 12542 13378 51986 13614
rect 52222 13378 52306 13614
rect 52542 13378 91986 13614
rect 92222 13378 92306 13614
rect 92542 13378 131986 13614
rect 132222 13378 132306 13614
rect 132542 13378 171986 13614
rect 172222 13378 172306 13614
rect 172542 13378 211986 13614
rect 212222 13378 212306 13614
rect 212542 13378 251986 13614
rect 252222 13378 252306 13614
rect 252542 13378 291986 13614
rect 292222 13378 292306 13614
rect 292542 13378 331986 13614
rect 332222 13378 332306 13614
rect 332542 13378 371986 13614
rect 372222 13378 372306 13614
rect 372542 13378 411986 13614
rect 412222 13378 412306 13614
rect 412542 13378 451986 13614
rect 452222 13378 452306 13614
rect 452542 13378 491986 13614
rect 492222 13378 492306 13614
rect 492542 13378 531986 13614
rect 532222 13378 532306 13614
rect 532542 13378 571986 13614
rect 572222 13378 572306 13614
rect 572542 13378 591102 13614
rect 591338 13378 591422 13614
rect 591658 13378 592650 13614
rect -8726 13294 592650 13378
rect -8726 13058 -7734 13294
rect -7498 13058 -7414 13294
rect -7178 13058 11986 13294
rect 12222 13058 12306 13294
rect 12542 13058 51986 13294
rect 52222 13058 52306 13294
rect 52542 13058 91986 13294
rect 92222 13058 92306 13294
rect 92542 13058 131986 13294
rect 132222 13058 132306 13294
rect 132542 13058 171986 13294
rect 172222 13058 172306 13294
rect 172542 13058 211986 13294
rect 212222 13058 212306 13294
rect 212542 13058 251986 13294
rect 252222 13058 252306 13294
rect 252542 13058 291986 13294
rect 292222 13058 292306 13294
rect 292542 13058 331986 13294
rect 332222 13058 332306 13294
rect 332542 13058 371986 13294
rect 372222 13058 372306 13294
rect 372542 13058 411986 13294
rect 412222 13058 412306 13294
rect 412542 13058 451986 13294
rect 452222 13058 452306 13294
rect 452542 13058 491986 13294
rect 492222 13058 492306 13294
rect 492542 13058 531986 13294
rect 532222 13058 532306 13294
rect 532542 13058 571986 13294
rect 572222 13058 572306 13294
rect 572542 13058 591102 13294
rect 591338 13058 591422 13294
rect 591658 13058 592650 13294
rect -8726 13026 592650 13058
rect -6806 9894 590730 9926
rect -6806 9658 -5814 9894
rect -5578 9658 -5494 9894
rect -5258 9658 8266 9894
rect 8502 9658 8586 9894
rect 8822 9658 48266 9894
rect 48502 9658 48586 9894
rect 48822 9658 88266 9894
rect 88502 9658 88586 9894
rect 88822 9658 128266 9894
rect 128502 9658 128586 9894
rect 128822 9658 168266 9894
rect 168502 9658 168586 9894
rect 168822 9658 208266 9894
rect 208502 9658 208586 9894
rect 208822 9658 248266 9894
rect 248502 9658 248586 9894
rect 248822 9658 288266 9894
rect 288502 9658 288586 9894
rect 288822 9658 328266 9894
rect 328502 9658 328586 9894
rect 328822 9658 368266 9894
rect 368502 9658 368586 9894
rect 368822 9658 408266 9894
rect 408502 9658 408586 9894
rect 408822 9658 448266 9894
rect 448502 9658 448586 9894
rect 448822 9658 488266 9894
rect 488502 9658 488586 9894
rect 488822 9658 528266 9894
rect 528502 9658 528586 9894
rect 528822 9658 568266 9894
rect 568502 9658 568586 9894
rect 568822 9658 589182 9894
rect 589418 9658 589502 9894
rect 589738 9658 590730 9894
rect -6806 9574 590730 9658
rect -6806 9338 -5814 9574
rect -5578 9338 -5494 9574
rect -5258 9338 8266 9574
rect 8502 9338 8586 9574
rect 8822 9338 48266 9574
rect 48502 9338 48586 9574
rect 48822 9338 88266 9574
rect 88502 9338 88586 9574
rect 88822 9338 128266 9574
rect 128502 9338 128586 9574
rect 128822 9338 168266 9574
rect 168502 9338 168586 9574
rect 168822 9338 208266 9574
rect 208502 9338 208586 9574
rect 208822 9338 248266 9574
rect 248502 9338 248586 9574
rect 248822 9338 288266 9574
rect 288502 9338 288586 9574
rect 288822 9338 328266 9574
rect 328502 9338 328586 9574
rect 328822 9338 368266 9574
rect 368502 9338 368586 9574
rect 368822 9338 408266 9574
rect 408502 9338 408586 9574
rect 408822 9338 448266 9574
rect 448502 9338 448586 9574
rect 448822 9338 488266 9574
rect 488502 9338 488586 9574
rect 488822 9338 528266 9574
rect 528502 9338 528586 9574
rect 528822 9338 568266 9574
rect 568502 9338 568586 9574
rect 568822 9338 589182 9574
rect 589418 9338 589502 9574
rect 589738 9338 590730 9574
rect -6806 9306 590730 9338
rect -4886 6174 588810 6206
rect -4886 5938 -3894 6174
rect -3658 5938 -3574 6174
rect -3338 5938 4546 6174
rect 4782 5938 4866 6174
rect 5102 5938 44546 6174
rect 44782 5938 44866 6174
rect 45102 5938 84546 6174
rect 84782 5938 84866 6174
rect 85102 5938 124546 6174
rect 124782 5938 124866 6174
rect 125102 5938 164546 6174
rect 164782 5938 164866 6174
rect 165102 5938 204546 6174
rect 204782 5938 204866 6174
rect 205102 5938 244546 6174
rect 244782 5938 244866 6174
rect 245102 5938 284546 6174
rect 284782 5938 284866 6174
rect 285102 5938 324546 6174
rect 324782 5938 324866 6174
rect 325102 5938 364546 6174
rect 364782 5938 364866 6174
rect 365102 5938 404546 6174
rect 404782 5938 404866 6174
rect 405102 5938 444546 6174
rect 444782 5938 444866 6174
rect 445102 5938 484546 6174
rect 484782 5938 484866 6174
rect 485102 5938 524546 6174
rect 524782 5938 524866 6174
rect 525102 5938 564546 6174
rect 564782 5938 564866 6174
rect 565102 5938 587262 6174
rect 587498 5938 587582 6174
rect 587818 5938 588810 6174
rect -4886 5854 588810 5938
rect -4886 5618 -3894 5854
rect -3658 5618 -3574 5854
rect -3338 5618 4546 5854
rect 4782 5618 4866 5854
rect 5102 5618 44546 5854
rect 44782 5618 44866 5854
rect 45102 5618 84546 5854
rect 84782 5618 84866 5854
rect 85102 5618 124546 5854
rect 124782 5618 124866 5854
rect 125102 5618 164546 5854
rect 164782 5618 164866 5854
rect 165102 5618 204546 5854
rect 204782 5618 204866 5854
rect 205102 5618 244546 5854
rect 244782 5618 244866 5854
rect 245102 5618 284546 5854
rect 284782 5618 284866 5854
rect 285102 5618 324546 5854
rect 324782 5618 324866 5854
rect 325102 5618 364546 5854
rect 364782 5618 364866 5854
rect 365102 5618 404546 5854
rect 404782 5618 404866 5854
rect 405102 5618 444546 5854
rect 444782 5618 444866 5854
rect 445102 5618 484546 5854
rect 484782 5618 484866 5854
rect 485102 5618 524546 5854
rect 524782 5618 524866 5854
rect 525102 5618 564546 5854
rect 564782 5618 564866 5854
rect 565102 5618 587262 5854
rect 587498 5618 587582 5854
rect 587818 5618 588810 5854
rect -4886 5586 588810 5618
rect -2966 2454 586890 2486
rect -2966 2218 -1974 2454
rect -1738 2218 -1654 2454
rect -1418 2218 826 2454
rect 1062 2218 1146 2454
rect 1382 2218 40826 2454
rect 41062 2218 41146 2454
rect 41382 2218 80826 2454
rect 81062 2218 81146 2454
rect 81382 2218 120826 2454
rect 121062 2218 121146 2454
rect 121382 2218 160826 2454
rect 161062 2218 161146 2454
rect 161382 2218 200826 2454
rect 201062 2218 201146 2454
rect 201382 2218 240826 2454
rect 241062 2218 241146 2454
rect 241382 2218 280826 2454
rect 281062 2218 281146 2454
rect 281382 2218 320826 2454
rect 321062 2218 321146 2454
rect 321382 2218 360826 2454
rect 361062 2218 361146 2454
rect 361382 2218 400826 2454
rect 401062 2218 401146 2454
rect 401382 2218 440826 2454
rect 441062 2218 441146 2454
rect 441382 2218 480826 2454
rect 481062 2218 481146 2454
rect 481382 2218 520826 2454
rect 521062 2218 521146 2454
rect 521382 2218 560826 2454
rect 561062 2218 561146 2454
rect 561382 2218 585342 2454
rect 585578 2218 585662 2454
rect 585898 2218 586890 2454
rect -2966 2134 586890 2218
rect -2966 1898 -1974 2134
rect -1738 1898 -1654 2134
rect -1418 1898 826 2134
rect 1062 1898 1146 2134
rect 1382 1898 40826 2134
rect 41062 1898 41146 2134
rect 41382 1898 80826 2134
rect 81062 1898 81146 2134
rect 81382 1898 120826 2134
rect 121062 1898 121146 2134
rect 121382 1898 160826 2134
rect 161062 1898 161146 2134
rect 161382 1898 200826 2134
rect 201062 1898 201146 2134
rect 201382 1898 240826 2134
rect 241062 1898 241146 2134
rect 241382 1898 280826 2134
rect 281062 1898 281146 2134
rect 281382 1898 320826 2134
rect 321062 1898 321146 2134
rect 321382 1898 360826 2134
rect 361062 1898 361146 2134
rect 361382 1898 400826 2134
rect 401062 1898 401146 2134
rect 401382 1898 440826 2134
rect 441062 1898 441146 2134
rect 441382 1898 480826 2134
rect 481062 1898 481146 2134
rect 481382 1898 520826 2134
rect 521062 1898 521146 2134
rect 521382 1898 560826 2134
rect 561062 1898 561146 2134
rect 561382 1898 585342 2134
rect 585578 1898 585662 2134
rect 585898 1898 586890 2134
rect -2966 1866 586890 1898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 826 -346
rect 1062 -582 1146 -346
rect 1382 -582 40826 -346
rect 41062 -582 41146 -346
rect 41382 -582 80826 -346
rect 81062 -582 81146 -346
rect 81382 -582 120826 -346
rect 121062 -582 121146 -346
rect 121382 -582 160826 -346
rect 161062 -582 161146 -346
rect 161382 -582 200826 -346
rect 201062 -582 201146 -346
rect 201382 -582 240826 -346
rect 241062 -582 241146 -346
rect 241382 -582 280826 -346
rect 281062 -582 281146 -346
rect 281382 -582 320826 -346
rect 321062 -582 321146 -346
rect 321382 -582 360826 -346
rect 361062 -582 361146 -346
rect 361382 -582 400826 -346
rect 401062 -582 401146 -346
rect 401382 -582 440826 -346
rect 441062 -582 441146 -346
rect 441382 -582 480826 -346
rect 481062 -582 481146 -346
rect 481382 -582 520826 -346
rect 521062 -582 521146 -346
rect 521382 -582 560826 -346
rect 561062 -582 561146 -346
rect 561382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 826 -666
rect 1062 -902 1146 -666
rect 1382 -902 40826 -666
rect 41062 -902 41146 -666
rect 41382 -902 80826 -666
rect 81062 -902 81146 -666
rect 81382 -902 120826 -666
rect 121062 -902 121146 -666
rect 121382 -902 160826 -666
rect 161062 -902 161146 -666
rect 161382 -902 200826 -666
rect 201062 -902 201146 -666
rect 201382 -902 240826 -666
rect 241062 -902 241146 -666
rect 241382 -902 280826 -666
rect 281062 -902 281146 -666
rect 281382 -902 320826 -666
rect 321062 -902 321146 -666
rect 321382 -902 360826 -666
rect 361062 -902 361146 -666
rect 361382 -902 400826 -666
rect 401062 -902 401146 -666
rect 401382 -902 440826 -666
rect 441062 -902 441146 -666
rect 441382 -902 480826 -666
rect 481062 -902 481146 -666
rect 481382 -902 520826 -666
rect 521062 -902 521146 -666
rect 521382 -902 560826 -666
rect 561062 -902 561146 -666
rect 561382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 20826 -1306
rect 21062 -1542 21146 -1306
rect 21382 -1542 60826 -1306
rect 61062 -1542 61146 -1306
rect 61382 -1542 100826 -1306
rect 101062 -1542 101146 -1306
rect 101382 -1542 140826 -1306
rect 141062 -1542 141146 -1306
rect 141382 -1542 180826 -1306
rect 181062 -1542 181146 -1306
rect 181382 -1542 220826 -1306
rect 221062 -1542 221146 -1306
rect 221382 -1542 260826 -1306
rect 261062 -1542 261146 -1306
rect 261382 -1542 300826 -1306
rect 301062 -1542 301146 -1306
rect 301382 -1542 340826 -1306
rect 341062 -1542 341146 -1306
rect 341382 -1542 380826 -1306
rect 381062 -1542 381146 -1306
rect 381382 -1542 420826 -1306
rect 421062 -1542 421146 -1306
rect 421382 -1542 460826 -1306
rect 461062 -1542 461146 -1306
rect 461382 -1542 500826 -1306
rect 501062 -1542 501146 -1306
rect 501382 -1542 540826 -1306
rect 541062 -1542 541146 -1306
rect 541382 -1542 580826 -1306
rect 581062 -1542 581146 -1306
rect 581382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 20826 -1626
rect 21062 -1862 21146 -1626
rect 21382 -1862 60826 -1626
rect 61062 -1862 61146 -1626
rect 61382 -1862 100826 -1626
rect 101062 -1862 101146 -1626
rect 101382 -1862 140826 -1626
rect 141062 -1862 141146 -1626
rect 141382 -1862 180826 -1626
rect 181062 -1862 181146 -1626
rect 181382 -1862 220826 -1626
rect 221062 -1862 221146 -1626
rect 221382 -1862 260826 -1626
rect 261062 -1862 261146 -1626
rect 261382 -1862 300826 -1626
rect 301062 -1862 301146 -1626
rect 301382 -1862 340826 -1626
rect 341062 -1862 341146 -1626
rect 341382 -1862 380826 -1626
rect 381062 -1862 381146 -1626
rect 381382 -1862 420826 -1626
rect 421062 -1862 421146 -1626
rect 421382 -1862 460826 -1626
rect 461062 -1862 461146 -1626
rect 461382 -1862 500826 -1626
rect 501062 -1862 501146 -1626
rect 501382 -1862 540826 -1626
rect 541062 -1862 541146 -1626
rect 541382 -1862 580826 -1626
rect 581062 -1862 581146 -1626
rect 581382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 4546 -2266
rect 4782 -2502 4866 -2266
rect 5102 -2502 44546 -2266
rect 44782 -2502 44866 -2266
rect 45102 -2502 84546 -2266
rect 84782 -2502 84866 -2266
rect 85102 -2502 124546 -2266
rect 124782 -2502 124866 -2266
rect 125102 -2502 164546 -2266
rect 164782 -2502 164866 -2266
rect 165102 -2502 204546 -2266
rect 204782 -2502 204866 -2266
rect 205102 -2502 244546 -2266
rect 244782 -2502 244866 -2266
rect 245102 -2502 284546 -2266
rect 284782 -2502 284866 -2266
rect 285102 -2502 324546 -2266
rect 324782 -2502 324866 -2266
rect 325102 -2502 364546 -2266
rect 364782 -2502 364866 -2266
rect 365102 -2502 404546 -2266
rect 404782 -2502 404866 -2266
rect 405102 -2502 444546 -2266
rect 444782 -2502 444866 -2266
rect 445102 -2502 484546 -2266
rect 484782 -2502 484866 -2266
rect 485102 -2502 524546 -2266
rect 524782 -2502 524866 -2266
rect 525102 -2502 564546 -2266
rect 564782 -2502 564866 -2266
rect 565102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 4546 -2586
rect 4782 -2822 4866 -2586
rect 5102 -2822 44546 -2586
rect 44782 -2822 44866 -2586
rect 45102 -2822 84546 -2586
rect 84782 -2822 84866 -2586
rect 85102 -2822 124546 -2586
rect 124782 -2822 124866 -2586
rect 125102 -2822 164546 -2586
rect 164782 -2822 164866 -2586
rect 165102 -2822 204546 -2586
rect 204782 -2822 204866 -2586
rect 205102 -2822 244546 -2586
rect 244782 -2822 244866 -2586
rect 245102 -2822 284546 -2586
rect 284782 -2822 284866 -2586
rect 285102 -2822 324546 -2586
rect 324782 -2822 324866 -2586
rect 325102 -2822 364546 -2586
rect 364782 -2822 364866 -2586
rect 365102 -2822 404546 -2586
rect 404782 -2822 404866 -2586
rect 405102 -2822 444546 -2586
rect 444782 -2822 444866 -2586
rect 445102 -2822 484546 -2586
rect 484782 -2822 484866 -2586
rect 485102 -2822 524546 -2586
rect 524782 -2822 524866 -2586
rect 525102 -2822 564546 -2586
rect 564782 -2822 564866 -2586
rect 565102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 24546 -3226
rect 24782 -3462 24866 -3226
rect 25102 -3462 64546 -3226
rect 64782 -3462 64866 -3226
rect 65102 -3462 104546 -3226
rect 104782 -3462 104866 -3226
rect 105102 -3462 144546 -3226
rect 144782 -3462 144866 -3226
rect 145102 -3462 184546 -3226
rect 184782 -3462 184866 -3226
rect 185102 -3462 224546 -3226
rect 224782 -3462 224866 -3226
rect 225102 -3462 264546 -3226
rect 264782 -3462 264866 -3226
rect 265102 -3462 304546 -3226
rect 304782 -3462 304866 -3226
rect 305102 -3462 344546 -3226
rect 344782 -3462 344866 -3226
rect 345102 -3462 384546 -3226
rect 384782 -3462 384866 -3226
rect 385102 -3462 424546 -3226
rect 424782 -3462 424866 -3226
rect 425102 -3462 464546 -3226
rect 464782 -3462 464866 -3226
rect 465102 -3462 504546 -3226
rect 504782 -3462 504866 -3226
rect 505102 -3462 544546 -3226
rect 544782 -3462 544866 -3226
rect 545102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 24546 -3546
rect 24782 -3782 24866 -3546
rect 25102 -3782 64546 -3546
rect 64782 -3782 64866 -3546
rect 65102 -3782 104546 -3546
rect 104782 -3782 104866 -3546
rect 105102 -3782 144546 -3546
rect 144782 -3782 144866 -3546
rect 145102 -3782 184546 -3546
rect 184782 -3782 184866 -3546
rect 185102 -3782 224546 -3546
rect 224782 -3782 224866 -3546
rect 225102 -3782 264546 -3546
rect 264782 -3782 264866 -3546
rect 265102 -3782 304546 -3546
rect 304782 -3782 304866 -3546
rect 305102 -3782 344546 -3546
rect 344782 -3782 344866 -3546
rect 345102 -3782 384546 -3546
rect 384782 -3782 384866 -3546
rect 385102 -3782 424546 -3546
rect 424782 -3782 424866 -3546
rect 425102 -3782 464546 -3546
rect 464782 -3782 464866 -3546
rect 465102 -3782 504546 -3546
rect 504782 -3782 504866 -3546
rect 505102 -3782 544546 -3546
rect 544782 -3782 544866 -3546
rect 545102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 8266 -4186
rect 8502 -4422 8586 -4186
rect 8822 -4422 48266 -4186
rect 48502 -4422 48586 -4186
rect 48822 -4422 88266 -4186
rect 88502 -4422 88586 -4186
rect 88822 -4422 128266 -4186
rect 128502 -4422 128586 -4186
rect 128822 -4422 168266 -4186
rect 168502 -4422 168586 -4186
rect 168822 -4422 208266 -4186
rect 208502 -4422 208586 -4186
rect 208822 -4422 248266 -4186
rect 248502 -4422 248586 -4186
rect 248822 -4422 288266 -4186
rect 288502 -4422 288586 -4186
rect 288822 -4422 328266 -4186
rect 328502 -4422 328586 -4186
rect 328822 -4422 368266 -4186
rect 368502 -4422 368586 -4186
rect 368822 -4422 408266 -4186
rect 408502 -4422 408586 -4186
rect 408822 -4422 448266 -4186
rect 448502 -4422 448586 -4186
rect 448822 -4422 488266 -4186
rect 488502 -4422 488586 -4186
rect 488822 -4422 528266 -4186
rect 528502 -4422 528586 -4186
rect 528822 -4422 568266 -4186
rect 568502 -4422 568586 -4186
rect 568822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 8266 -4506
rect 8502 -4742 8586 -4506
rect 8822 -4742 48266 -4506
rect 48502 -4742 48586 -4506
rect 48822 -4742 88266 -4506
rect 88502 -4742 88586 -4506
rect 88822 -4742 128266 -4506
rect 128502 -4742 128586 -4506
rect 128822 -4742 168266 -4506
rect 168502 -4742 168586 -4506
rect 168822 -4742 208266 -4506
rect 208502 -4742 208586 -4506
rect 208822 -4742 248266 -4506
rect 248502 -4742 248586 -4506
rect 248822 -4742 288266 -4506
rect 288502 -4742 288586 -4506
rect 288822 -4742 328266 -4506
rect 328502 -4742 328586 -4506
rect 328822 -4742 368266 -4506
rect 368502 -4742 368586 -4506
rect 368822 -4742 408266 -4506
rect 408502 -4742 408586 -4506
rect 408822 -4742 448266 -4506
rect 448502 -4742 448586 -4506
rect 448822 -4742 488266 -4506
rect 488502 -4742 488586 -4506
rect 488822 -4742 528266 -4506
rect 528502 -4742 528586 -4506
rect 528822 -4742 568266 -4506
rect 568502 -4742 568586 -4506
rect 568822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 28266 -5146
rect 28502 -5382 28586 -5146
rect 28822 -5382 68266 -5146
rect 68502 -5382 68586 -5146
rect 68822 -5382 108266 -5146
rect 108502 -5382 108586 -5146
rect 108822 -5382 148266 -5146
rect 148502 -5382 148586 -5146
rect 148822 -5382 188266 -5146
rect 188502 -5382 188586 -5146
rect 188822 -5382 228266 -5146
rect 228502 -5382 228586 -5146
rect 228822 -5382 268266 -5146
rect 268502 -5382 268586 -5146
rect 268822 -5382 308266 -5146
rect 308502 -5382 308586 -5146
rect 308822 -5382 348266 -5146
rect 348502 -5382 348586 -5146
rect 348822 -5382 388266 -5146
rect 388502 -5382 388586 -5146
rect 388822 -5382 428266 -5146
rect 428502 -5382 428586 -5146
rect 428822 -5382 468266 -5146
rect 468502 -5382 468586 -5146
rect 468822 -5382 508266 -5146
rect 508502 -5382 508586 -5146
rect 508822 -5382 548266 -5146
rect 548502 -5382 548586 -5146
rect 548822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 28266 -5466
rect 28502 -5702 28586 -5466
rect 28822 -5702 68266 -5466
rect 68502 -5702 68586 -5466
rect 68822 -5702 108266 -5466
rect 108502 -5702 108586 -5466
rect 108822 -5702 148266 -5466
rect 148502 -5702 148586 -5466
rect 148822 -5702 188266 -5466
rect 188502 -5702 188586 -5466
rect 188822 -5702 228266 -5466
rect 228502 -5702 228586 -5466
rect 228822 -5702 268266 -5466
rect 268502 -5702 268586 -5466
rect 268822 -5702 308266 -5466
rect 308502 -5702 308586 -5466
rect 308822 -5702 348266 -5466
rect 348502 -5702 348586 -5466
rect 348822 -5702 388266 -5466
rect 388502 -5702 388586 -5466
rect 388822 -5702 428266 -5466
rect 428502 -5702 428586 -5466
rect 428822 -5702 468266 -5466
rect 468502 -5702 468586 -5466
rect 468822 -5702 508266 -5466
rect 508502 -5702 508586 -5466
rect 508822 -5702 548266 -5466
rect 548502 -5702 548586 -5466
rect 548822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 11986 -6106
rect 12222 -6342 12306 -6106
rect 12542 -6342 51986 -6106
rect 52222 -6342 52306 -6106
rect 52542 -6342 91986 -6106
rect 92222 -6342 92306 -6106
rect 92542 -6342 131986 -6106
rect 132222 -6342 132306 -6106
rect 132542 -6342 171986 -6106
rect 172222 -6342 172306 -6106
rect 172542 -6342 211986 -6106
rect 212222 -6342 212306 -6106
rect 212542 -6342 251986 -6106
rect 252222 -6342 252306 -6106
rect 252542 -6342 291986 -6106
rect 292222 -6342 292306 -6106
rect 292542 -6342 331986 -6106
rect 332222 -6342 332306 -6106
rect 332542 -6342 371986 -6106
rect 372222 -6342 372306 -6106
rect 372542 -6342 411986 -6106
rect 412222 -6342 412306 -6106
rect 412542 -6342 451986 -6106
rect 452222 -6342 452306 -6106
rect 452542 -6342 491986 -6106
rect 492222 -6342 492306 -6106
rect 492542 -6342 531986 -6106
rect 532222 -6342 532306 -6106
rect 532542 -6342 571986 -6106
rect 572222 -6342 572306 -6106
rect 572542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 11986 -6426
rect 12222 -6662 12306 -6426
rect 12542 -6662 51986 -6426
rect 52222 -6662 52306 -6426
rect 52542 -6662 91986 -6426
rect 92222 -6662 92306 -6426
rect 92542 -6662 131986 -6426
rect 132222 -6662 132306 -6426
rect 132542 -6662 171986 -6426
rect 172222 -6662 172306 -6426
rect 172542 -6662 211986 -6426
rect 212222 -6662 212306 -6426
rect 212542 -6662 251986 -6426
rect 252222 -6662 252306 -6426
rect 252542 -6662 291986 -6426
rect 292222 -6662 292306 -6426
rect 292542 -6662 331986 -6426
rect 332222 -6662 332306 -6426
rect 332542 -6662 371986 -6426
rect 372222 -6662 372306 -6426
rect 372542 -6662 411986 -6426
rect 412222 -6662 412306 -6426
rect 412542 -6662 451986 -6426
rect 452222 -6662 452306 -6426
rect 452542 -6662 491986 -6426
rect 492222 -6662 492306 -6426
rect 492542 -6662 531986 -6426
rect 532222 -6662 532306 -6426
rect 532542 -6662 571986 -6426
rect 572222 -6662 572306 -6426
rect 572542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 31986 -7066
rect 32222 -7302 32306 -7066
rect 32542 -7302 71986 -7066
rect 72222 -7302 72306 -7066
rect 72542 -7302 111986 -7066
rect 112222 -7302 112306 -7066
rect 112542 -7302 151986 -7066
rect 152222 -7302 152306 -7066
rect 152542 -7302 191986 -7066
rect 192222 -7302 192306 -7066
rect 192542 -7302 231986 -7066
rect 232222 -7302 232306 -7066
rect 232542 -7302 271986 -7066
rect 272222 -7302 272306 -7066
rect 272542 -7302 311986 -7066
rect 312222 -7302 312306 -7066
rect 312542 -7302 351986 -7066
rect 352222 -7302 352306 -7066
rect 352542 -7302 391986 -7066
rect 392222 -7302 392306 -7066
rect 392542 -7302 431986 -7066
rect 432222 -7302 432306 -7066
rect 432542 -7302 471986 -7066
rect 472222 -7302 472306 -7066
rect 472542 -7302 511986 -7066
rect 512222 -7302 512306 -7066
rect 512542 -7302 551986 -7066
rect 552222 -7302 552306 -7066
rect 552542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 31986 -7386
rect 32222 -7622 32306 -7386
rect 32542 -7622 71986 -7386
rect 72222 -7622 72306 -7386
rect 72542 -7622 111986 -7386
rect 112222 -7622 112306 -7386
rect 112542 -7622 151986 -7386
rect 152222 -7622 152306 -7386
rect 152542 -7622 191986 -7386
rect 192222 -7622 192306 -7386
rect 192542 -7622 231986 -7386
rect 232222 -7622 232306 -7386
rect 232542 -7622 271986 -7386
rect 272222 -7622 272306 -7386
rect 272542 -7622 311986 -7386
rect 312222 -7622 312306 -7386
rect 312542 -7622 351986 -7386
rect 352222 -7622 352306 -7386
rect 352542 -7622 391986 -7386
rect 392222 -7622 392306 -7386
rect 392542 -7622 431986 -7386
rect 432222 -7622 432306 -7386
rect 432542 -7622 471986 -7386
rect 472222 -7622 472306 -7386
rect 472542 -7622 511986 -7386
rect 512222 -7622 512306 -7386
rect 512542 -7622 551986 -7386
rect 552222 -7622 552306 -7386
rect 552542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use multiplier  MULT
timestamp 1641153771
transform 1 0 120000 0 1 120000
box 0 0 200000 200000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 1866 586890 2486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 41866 586890 42486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 81866 586890 82486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 121866 586890 122486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 161866 586890 162486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 201866 586890 202486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 241866 586890 242486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 281866 586890 282486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 321866 586890 322486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 361866 586890 362486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 401866 586890 402486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 441866 586890 442486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 481866 586890 482486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 521866 586890 522486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 561866 586890 562486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 601866 586890 602486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 641866 586890 642486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 681866 586890 682486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 794 -1894 1414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 40794 -1894 41414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 80794 -1894 81414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 120794 -1894 121414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 160794 -1894 161414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 200794 -1894 201414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 240794 -1894 241414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 280794 -1894 281414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 320794 -1894 321414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 360794 -1894 361414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 400794 -1894 401414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 440794 -1894 441414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 480794 -1894 481414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 520794 -1894 521414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 560794 -1894 561414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 5586 588810 6206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 45586 588810 46206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 85586 588810 86206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 125586 588810 126206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 165586 588810 166206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 205586 588810 206206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 245586 588810 246206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 285586 588810 286206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 325586 588810 326206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 365586 588810 366206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 405586 588810 406206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 445586 588810 446206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 485586 588810 486206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 525586 588810 526206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 565586 588810 566206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 605586 588810 606206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 645586 588810 646206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 685586 588810 686206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 4514 -3814 5134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 44514 -3814 45134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 84514 -3814 85134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 124514 -3814 125134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 164514 -3814 165134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 204514 -3814 205134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 244514 -3814 245134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 284514 -3814 285134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 324514 -3814 325134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 364514 -3814 365134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 404514 -3814 405134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 444514 -3814 445134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 484514 -3814 485134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 524514 -3814 525134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 564514 -3814 565134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 9306 590730 9926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 49306 590730 49926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 89306 590730 89926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 129306 590730 129926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 169306 590730 169926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 209306 590730 209926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 249306 590730 249926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 289306 590730 289926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 329306 590730 329926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 369306 590730 369926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 409306 590730 409926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 449306 590730 449926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 489306 590730 489926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 529306 590730 529926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 569306 590730 569926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 609306 590730 609926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 649306 590730 649926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 689306 590730 689926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 8234 -5734 8854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 48234 -5734 48854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 88234 -5734 88854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 128234 -5734 128854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 168234 -5734 168854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 208234 -5734 208854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 248234 -5734 248854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 288234 -5734 288854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 328234 -5734 328854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 368234 -5734 368854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 408234 -5734 408854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 448234 -5734 448854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 488234 -5734 488854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 528234 -5734 528854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 568234 -5734 568854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 13026 592650 13646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 53026 592650 53646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 93026 592650 93646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 133026 592650 133646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 173026 592650 173646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 213026 592650 213646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 253026 592650 253646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 293026 592650 293646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 333026 592650 333646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 373026 592650 373646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 413026 592650 413646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 453026 592650 453646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 493026 592650 493646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 533026 592650 533646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 573026 592650 573646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 613026 592650 613646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 653026 592650 653646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 693026 592650 693646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 11954 -7654 12574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 51954 -7654 52574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 91954 -7654 92574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 131954 -7654 132574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 171954 -7654 172574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 211954 -7654 212574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 251954 -7654 252574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 291954 -7654 292574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 331954 -7654 332574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 371954 -7654 372574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 411954 -7654 412574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 451954 -7654 452574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 491954 -7654 492574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 531954 -7654 532574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 571954 -7654 572574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 29306 590730 29926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 69306 590730 69926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 109306 590730 109926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 149306 590730 149926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 189306 590730 189926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 229306 590730 229926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 269306 590730 269926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 309306 590730 309926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 349306 590730 349926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 389306 590730 389926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 429306 590730 429926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 469306 590730 469926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 509306 590730 509926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 549306 590730 549926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 589306 590730 589926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 629306 590730 629926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 669306 590730 669926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 28234 -5734 28854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 68234 -5734 68854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 108234 -5734 108854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 148234 -5734 148854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 188234 -5734 188854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 228234 -5734 228854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 268234 -5734 268854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 308234 -5734 308854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 348234 -5734 348854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 388234 -5734 388854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 428234 -5734 428854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 468234 -5734 468854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 508234 -5734 508854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 548234 -5734 548854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 33026 592650 33646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 73026 592650 73646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 113026 592650 113646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 153026 592650 153646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 193026 592650 193646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 233026 592650 233646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 273026 592650 273646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 313026 592650 313646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 353026 592650 353646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 393026 592650 393646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 433026 592650 433646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 473026 592650 473646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 513026 592650 513646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 553026 592650 553646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 593026 592650 593646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 633026 592650 633646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 673026 592650 673646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 31954 -7654 32574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 71954 -7654 72574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 111954 -7654 112574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 151954 -7654 152574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 191954 -7654 192574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 231954 -7654 232574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 271954 -7654 272574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 311954 -7654 312574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 351954 -7654 352574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 391954 -7654 392574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 431954 -7654 432574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 471954 -7654 472574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 511954 -7654 512574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 551954 -7654 552574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 21866 586890 22486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 61866 586890 62486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 101866 586890 102486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 141866 586890 142486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 181866 586890 182486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 221866 586890 222486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 261866 586890 262486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 301866 586890 302486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 341866 586890 342486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 381866 586890 382486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 421866 586890 422486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 461866 586890 462486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 501866 586890 502486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 541866 586890 542486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 581866 586890 582486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 621866 586890 622486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 661866 586890 662486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 20794 -1894 21414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 60794 -1894 61414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 100794 -1894 101414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 140794 -1894 141414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 180794 -1894 181414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 220794 -1894 221414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 260794 -1894 261414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 300794 -1894 301414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 340794 -1894 341414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 380794 -1894 381414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 420794 -1894 421414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 460794 -1894 461414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 500794 -1894 501414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 540794 -1894 541414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 580794 -1894 581414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 25586 588810 26206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 65586 588810 66206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 105586 588810 106206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 145586 588810 146206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 185586 588810 186206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 225586 588810 226206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 265586 588810 266206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 305586 588810 306206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 345586 588810 346206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 385586 588810 386206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 425586 588810 426206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 465586 588810 466206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 505586 588810 506206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 545586 588810 546206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 585586 588810 586206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 625586 588810 626206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 665586 588810 666206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 24514 -3814 25134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 64514 -3814 65134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 104514 -3814 105134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 144514 -3814 145134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 184514 -3814 185134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 224514 -3814 225134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 264514 -3814 265134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 304514 -3814 305134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 344514 -3814 345134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 384514 -3814 385134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 424514 -3814 425134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 464514 -3814 465134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 504514 -3814 505134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 544514 -3814 545134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
